VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 450.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 10.640 75.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 10.640 125.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 10.640 175.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 10.640 225.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 10.640 275.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 438.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 444.600 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.030 444.600 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 130.030 444.600 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 180.030 444.600 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 230.030 444.600 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 280.030 444.600 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 330.030 444.600 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 444.600 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 430.030 444.600 431.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 438.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 444.600 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 444.600 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 126.730 444.600 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 176.730 444.600 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 226.730 444.600 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 276.730 444.600 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.730 444.600 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 444.600 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 426.730 444.600 428.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 312.840 450.000 313.440 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 176.840 450.000 177.440 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 190.440 450.000 191.040 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 204.040 450.000 204.640 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 217.640 450.000 218.240 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 231.240 450.000 231.840 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 244.840 450.000 245.440 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 258.440 450.000 259.040 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 272.040 450.000 272.640 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 285.640 450.000 286.240 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 299.240 450.000 299.840 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 326.440 450.000 327.040 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 40.840 450.000 41.440 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 54.440 450.000 55.040 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 68.040 450.000 68.640 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 81.640 450.000 82.240 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 95.240 450.000 95.840 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 108.840 450.000 109.440 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 122.440 450.000 123.040 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 136.040 450.000 136.640 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 149.640 450.000 150.240 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 163.240 450.000 163.840 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 340.040 450.000 340.640 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 13.640 450.000 14.240 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 27.240 450.000 27.840 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.870 446.000 342.150 450.000 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 355.670 446.000 355.950 450.000 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 369.470 446.000 369.750 450.000 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 446.000 383.550 450.000 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 397.070 446.000 397.350 450.000 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 410.870 446.000 411.150 450.000 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 424.670 446.000 424.950 450.000 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 438.470 446.000 438.750 450.000 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 353.640 450.000 354.240 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 203.870 446.000 204.150 450.000 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 217.670 446.000 217.950 450.000 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 231.470 446.000 231.750 450.000 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 245.270 446.000 245.550 450.000 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 259.070 446.000 259.350 450.000 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 272.870 446.000 273.150 450.000 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 446.000 286.950 450.000 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 300.470 446.000 300.750 450.000 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 314.270 446.000 314.550 450.000 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 328.070 446.000 328.350 450.000 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 367.240 450.000 367.840 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 446.000 66.150 450.000 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.670 446.000 79.950 450.000 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 446.000 93.750 450.000 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 446.000 107.550 450.000 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 446.000 121.350 450.000 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.870 446.000 135.150 450.000 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.670 446.000 148.950 450.000 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.470 446.000 162.750 450.000 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 446.000 176.550 450.000 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 446.000 190.350 450.000 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 380.840 450.000 381.440 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 10.670 446.000 10.950 450.000 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 446.000 24.750 450.000 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 446.000 38.550 450.000 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.070 446.000 52.350 450.000 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 394.440 450.000 395.040 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 408.040 450.000 408.640 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 421.640 450.000 422.240 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 435.240 450.000 435.840 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 444.550 438.110 ;
      LAYER li1 ;
        RECT 5.520 10.795 444.360 438.005 ;
      LAYER met1 ;
        RECT 4.210 10.240 444.660 438.560 ;
      LAYER met2 ;
        RECT 4.230 445.720 10.390 446.490 ;
        RECT 11.230 445.720 24.190 446.490 ;
        RECT 25.030 445.720 37.990 446.490 ;
        RECT 38.830 445.720 51.790 446.490 ;
        RECT 52.630 445.720 65.590 446.490 ;
        RECT 66.430 445.720 79.390 446.490 ;
        RECT 80.230 445.720 93.190 446.490 ;
        RECT 94.030 445.720 106.990 446.490 ;
        RECT 107.830 445.720 120.790 446.490 ;
        RECT 121.630 445.720 134.590 446.490 ;
        RECT 135.430 445.720 148.390 446.490 ;
        RECT 149.230 445.720 162.190 446.490 ;
        RECT 163.030 445.720 175.990 446.490 ;
        RECT 176.830 445.720 189.790 446.490 ;
        RECT 190.630 445.720 203.590 446.490 ;
        RECT 204.430 445.720 217.390 446.490 ;
        RECT 218.230 445.720 231.190 446.490 ;
        RECT 232.030 445.720 244.990 446.490 ;
        RECT 245.830 445.720 258.790 446.490 ;
        RECT 259.630 445.720 272.590 446.490 ;
        RECT 273.430 445.720 286.390 446.490 ;
        RECT 287.230 445.720 300.190 446.490 ;
        RECT 301.030 445.720 313.990 446.490 ;
        RECT 314.830 445.720 327.790 446.490 ;
        RECT 328.630 445.720 341.590 446.490 ;
        RECT 342.430 445.720 355.390 446.490 ;
        RECT 356.230 445.720 369.190 446.490 ;
        RECT 370.030 445.720 382.990 446.490 ;
        RECT 383.830 445.720 396.790 446.490 ;
        RECT 397.630 445.720 410.590 446.490 ;
        RECT 411.430 445.720 424.390 446.490 ;
        RECT 425.230 445.720 438.190 446.490 ;
        RECT 439.030 445.720 444.260 446.490 ;
        RECT 4.230 4.280 444.260 445.720 ;
        RECT 4.230 3.670 10.850 4.280 ;
        RECT 11.690 3.670 24.190 4.280 ;
        RECT 25.030 3.670 37.530 4.280 ;
        RECT 38.370 3.670 50.870 4.280 ;
        RECT 51.710 3.670 64.210 4.280 ;
        RECT 65.050 3.670 77.550 4.280 ;
        RECT 78.390 3.670 90.890 4.280 ;
        RECT 91.730 3.670 104.230 4.280 ;
        RECT 105.070 3.670 117.570 4.280 ;
        RECT 118.410 3.670 130.910 4.280 ;
        RECT 131.750 3.670 144.250 4.280 ;
        RECT 145.090 3.670 157.590 4.280 ;
        RECT 158.430 3.670 170.930 4.280 ;
        RECT 171.770 3.670 184.270 4.280 ;
        RECT 185.110 3.670 197.610 4.280 ;
        RECT 198.450 3.670 210.950 4.280 ;
        RECT 211.790 3.670 224.290 4.280 ;
        RECT 225.130 3.670 237.630 4.280 ;
        RECT 238.470 3.670 250.970 4.280 ;
        RECT 251.810 3.670 264.310 4.280 ;
        RECT 265.150 3.670 277.650 4.280 ;
        RECT 278.490 3.670 290.990 4.280 ;
        RECT 291.830 3.670 304.330 4.280 ;
        RECT 305.170 3.670 317.670 4.280 ;
        RECT 318.510 3.670 331.010 4.280 ;
        RECT 331.850 3.670 344.350 4.280 ;
        RECT 345.190 3.670 357.690 4.280 ;
        RECT 358.530 3.670 371.030 4.280 ;
        RECT 371.870 3.670 384.370 4.280 ;
        RECT 385.210 3.670 397.710 4.280 ;
        RECT 398.550 3.670 411.050 4.280 ;
        RECT 411.890 3.670 424.390 4.280 ;
        RECT 425.230 3.670 437.730 4.280 ;
        RECT 438.570 3.670 444.260 4.280 ;
      LAYER met3 ;
        RECT 4.400 441.640 446.000 442.490 ;
        RECT 3.990 436.240 446.000 441.640 ;
        RECT 3.990 434.840 445.600 436.240 ;
        RECT 3.990 429.440 446.000 434.840 ;
        RECT 4.400 428.040 446.000 429.440 ;
        RECT 3.990 422.640 446.000 428.040 ;
        RECT 3.990 421.240 445.600 422.640 ;
        RECT 3.990 415.840 446.000 421.240 ;
        RECT 4.400 414.440 446.000 415.840 ;
        RECT 3.990 409.040 446.000 414.440 ;
        RECT 3.990 407.640 445.600 409.040 ;
        RECT 3.990 402.240 446.000 407.640 ;
        RECT 4.400 400.840 446.000 402.240 ;
        RECT 3.990 395.440 446.000 400.840 ;
        RECT 3.990 394.040 445.600 395.440 ;
        RECT 3.990 388.640 446.000 394.040 ;
        RECT 4.400 387.240 446.000 388.640 ;
        RECT 3.990 381.840 446.000 387.240 ;
        RECT 3.990 380.440 445.600 381.840 ;
        RECT 3.990 375.040 446.000 380.440 ;
        RECT 4.400 373.640 446.000 375.040 ;
        RECT 3.990 368.240 446.000 373.640 ;
        RECT 3.990 366.840 445.600 368.240 ;
        RECT 3.990 361.440 446.000 366.840 ;
        RECT 4.400 360.040 446.000 361.440 ;
        RECT 3.990 354.640 446.000 360.040 ;
        RECT 3.990 353.240 445.600 354.640 ;
        RECT 3.990 347.840 446.000 353.240 ;
        RECT 4.400 346.440 446.000 347.840 ;
        RECT 3.990 341.040 446.000 346.440 ;
        RECT 3.990 339.640 445.600 341.040 ;
        RECT 3.990 334.240 446.000 339.640 ;
        RECT 4.400 332.840 446.000 334.240 ;
        RECT 3.990 327.440 446.000 332.840 ;
        RECT 3.990 326.040 445.600 327.440 ;
        RECT 3.990 320.640 446.000 326.040 ;
        RECT 4.400 319.240 446.000 320.640 ;
        RECT 3.990 313.840 446.000 319.240 ;
        RECT 3.990 312.440 445.600 313.840 ;
        RECT 3.990 307.040 446.000 312.440 ;
        RECT 4.400 305.640 446.000 307.040 ;
        RECT 3.990 300.240 446.000 305.640 ;
        RECT 3.990 298.840 445.600 300.240 ;
        RECT 3.990 293.440 446.000 298.840 ;
        RECT 4.400 292.040 446.000 293.440 ;
        RECT 3.990 286.640 446.000 292.040 ;
        RECT 3.990 285.240 445.600 286.640 ;
        RECT 3.990 279.840 446.000 285.240 ;
        RECT 4.400 278.440 446.000 279.840 ;
        RECT 3.990 273.040 446.000 278.440 ;
        RECT 3.990 271.640 445.600 273.040 ;
        RECT 3.990 266.240 446.000 271.640 ;
        RECT 4.400 264.840 446.000 266.240 ;
        RECT 3.990 259.440 446.000 264.840 ;
        RECT 3.990 258.040 445.600 259.440 ;
        RECT 3.990 252.640 446.000 258.040 ;
        RECT 4.400 251.240 446.000 252.640 ;
        RECT 3.990 245.840 446.000 251.240 ;
        RECT 3.990 244.440 445.600 245.840 ;
        RECT 3.990 239.040 446.000 244.440 ;
        RECT 4.400 237.640 446.000 239.040 ;
        RECT 3.990 232.240 446.000 237.640 ;
        RECT 3.990 230.840 445.600 232.240 ;
        RECT 3.990 225.440 446.000 230.840 ;
        RECT 4.400 224.040 446.000 225.440 ;
        RECT 3.990 218.640 446.000 224.040 ;
        RECT 3.990 217.240 445.600 218.640 ;
        RECT 3.990 211.840 446.000 217.240 ;
        RECT 4.400 210.440 446.000 211.840 ;
        RECT 3.990 205.040 446.000 210.440 ;
        RECT 3.990 203.640 445.600 205.040 ;
        RECT 3.990 198.240 446.000 203.640 ;
        RECT 4.400 196.840 446.000 198.240 ;
        RECT 3.990 191.440 446.000 196.840 ;
        RECT 3.990 190.040 445.600 191.440 ;
        RECT 3.990 184.640 446.000 190.040 ;
        RECT 4.400 183.240 446.000 184.640 ;
        RECT 3.990 177.840 446.000 183.240 ;
        RECT 3.990 176.440 445.600 177.840 ;
        RECT 3.990 171.040 446.000 176.440 ;
        RECT 4.400 169.640 446.000 171.040 ;
        RECT 3.990 164.240 446.000 169.640 ;
        RECT 3.990 162.840 445.600 164.240 ;
        RECT 3.990 157.440 446.000 162.840 ;
        RECT 4.400 156.040 446.000 157.440 ;
        RECT 3.990 150.640 446.000 156.040 ;
        RECT 3.990 149.240 445.600 150.640 ;
        RECT 3.990 143.840 446.000 149.240 ;
        RECT 4.400 142.440 446.000 143.840 ;
        RECT 3.990 137.040 446.000 142.440 ;
        RECT 3.990 135.640 445.600 137.040 ;
        RECT 3.990 130.240 446.000 135.640 ;
        RECT 4.400 128.840 446.000 130.240 ;
        RECT 3.990 123.440 446.000 128.840 ;
        RECT 3.990 122.040 445.600 123.440 ;
        RECT 3.990 116.640 446.000 122.040 ;
        RECT 4.400 115.240 446.000 116.640 ;
        RECT 3.990 109.840 446.000 115.240 ;
        RECT 3.990 108.440 445.600 109.840 ;
        RECT 3.990 103.040 446.000 108.440 ;
        RECT 4.400 101.640 446.000 103.040 ;
        RECT 3.990 96.240 446.000 101.640 ;
        RECT 3.990 94.840 445.600 96.240 ;
        RECT 3.990 89.440 446.000 94.840 ;
        RECT 4.400 88.040 446.000 89.440 ;
        RECT 3.990 82.640 446.000 88.040 ;
        RECT 3.990 81.240 445.600 82.640 ;
        RECT 3.990 75.840 446.000 81.240 ;
        RECT 4.400 74.440 446.000 75.840 ;
        RECT 3.990 69.040 446.000 74.440 ;
        RECT 3.990 67.640 445.600 69.040 ;
        RECT 3.990 62.240 446.000 67.640 ;
        RECT 4.400 60.840 446.000 62.240 ;
        RECT 3.990 55.440 446.000 60.840 ;
        RECT 3.990 54.040 445.600 55.440 ;
        RECT 3.990 48.640 446.000 54.040 ;
        RECT 4.400 47.240 446.000 48.640 ;
        RECT 3.990 41.840 446.000 47.240 ;
        RECT 3.990 40.440 445.600 41.840 ;
        RECT 3.990 35.040 446.000 40.440 ;
        RECT 4.400 33.640 446.000 35.040 ;
        RECT 3.990 28.240 446.000 33.640 ;
        RECT 3.990 26.840 445.600 28.240 ;
        RECT 3.990 21.440 446.000 26.840 ;
        RECT 4.400 20.040 446.000 21.440 ;
        RECT 3.990 14.640 446.000 20.040 ;
        RECT 3.990 13.240 445.600 14.640 ;
        RECT 3.990 7.840 446.000 13.240 ;
        RECT 4.400 6.990 446.000 7.840 ;
      LAYER met4 ;
        RECT 15.935 13.775 20.640 417.345 ;
        RECT 23.040 13.775 23.940 417.345 ;
        RECT 26.340 13.775 70.640 417.345 ;
        RECT 73.040 13.775 73.940 417.345 ;
        RECT 76.340 13.775 120.640 417.345 ;
        RECT 123.040 13.775 123.940 417.345 ;
        RECT 126.340 13.775 170.640 417.345 ;
        RECT 173.040 13.775 173.940 417.345 ;
        RECT 176.340 13.775 220.640 417.345 ;
        RECT 223.040 13.775 223.940 417.345 ;
        RECT 226.340 13.775 270.640 417.345 ;
        RECT 273.040 13.775 273.940 417.345 ;
        RECT 276.340 13.775 320.640 417.345 ;
        RECT 323.040 13.775 323.940 417.345 ;
        RECT 326.340 13.775 370.640 417.345 ;
        RECT 373.040 13.775 373.940 417.345 ;
        RECT 376.340 13.775 420.640 417.345 ;
        RECT 423.040 13.775 423.940 417.345 ;
        RECT 426.340 13.775 430.265 417.345 ;
  END
END pipelined_mult
END LIBRARY

