VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mult_16x16
  CLASS BLOCK ;
  FOREIGN mult_16x16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 225.000 BY 225.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 212.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 219.660 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 219.660 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 212.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 212.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 219.660 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 219.660 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 199.730 221.000 200.010 225.000 ;
    END
  END clk
  PIN in1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 221.000 29.350 225.000 ;
    END
  END in1[0]
  PIN in1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END in1[10]
  PIN in1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END in1[11]
  PIN in1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END in1[12]
  PIN in1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END in1[13]
  PIN in1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END in1[14]
  PIN in1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END in1[15]
  PIN in1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 221.000 39.010 225.000 ;
    END
  END in1[1]
  PIN in1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 221.000 45.450 225.000 ;
    END
  END in1[2]
  PIN in1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 221.000 51.890 225.000 ;
    END
  END in1[3]
  PIN in1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.590 221.000 80.870 225.000 ;
    END
  END in1[4]
  PIN in1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 221.000 103.410 225.000 ;
    END
  END in1[5]
  PIN in1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 221.000 125.840 225.000 126.440 ;
    END
  END in1[6]
  PIN in1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.090 221.000 161.370 225.000 ;
    END
  END in1[7]
  PIN in1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 221.000 119.040 225.000 119.640 ;
    END
  END in1[8]
  PIN in1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END in1[9]
  PIN in2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 221.000 129.240 225.000 129.840 ;
    END
  END in2[0]
  PIN in2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END in2[10]
  PIN in2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END in2[11]
  PIN in2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END in2[12]
  PIN in2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END in2[13]
  PIN in2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END in2[14]
  PIN in2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END in2[15]
  PIN in2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 221.000 136.040 225.000 136.640 ;
    END
  END in2[1]
  PIN in2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 221.000 139.440 225.000 140.040 ;
    END
  END in2[2]
  PIN in2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.790 221.000 113.070 225.000 ;
    END
  END in2[3]
  PIN in2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 221.000 90.530 225.000 ;
    END
  END in2[4]
  PIN in2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 221.000 116.290 225.000 ;
    END
  END in2[5]
  PIN in2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.030 221.000 87.310 225.000 ;
    END
  END in2[6]
  PIN in2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.470 221.000 93.750 225.000 ;
    END
  END in2[7]
  PIN in2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 221.000 84.090 225.000 ;
    END
  END in2[8]
  PIN in2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 221.000 32.570 225.000 ;
    END
  END in2[9]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 142.840 225.000 143.440 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 221.000 119.510 225.000 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 221.000 58.330 225.000 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 221.000 48.670 225.000 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 221.000 35.790 225.000 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 153.040 225.000 153.640 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 149.640 225.000 150.240 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END out[31]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 159.840 225.000 160.440 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 173.440 225.000 174.040 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 187.040 225.000 187.640 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 197.240 225.000 197.840 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 221.000 204.040 225.000 204.640 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 221.000 203.230 225.000 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 221.000 132.390 225.000 ;
    END
  END out[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 221.000 206.450 225.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 219.610 212.245 ;
      LAYER li1 ;
        RECT 5.520 10.795 219.420 212.245 ;
      LAYER met1 ;
        RECT 4.210 10.640 219.420 213.820 ;
      LAYER met2 ;
        RECT 4.230 220.720 28.790 221.525 ;
        RECT 29.630 220.720 32.010 221.525 ;
        RECT 32.850 220.720 35.230 221.525 ;
        RECT 36.070 220.720 38.450 221.525 ;
        RECT 39.290 220.720 44.890 221.525 ;
        RECT 45.730 220.720 48.110 221.525 ;
        RECT 48.950 220.720 51.330 221.525 ;
        RECT 52.170 220.720 57.770 221.525 ;
        RECT 58.610 220.720 80.310 221.525 ;
        RECT 81.150 220.720 83.530 221.525 ;
        RECT 84.370 220.720 86.750 221.525 ;
        RECT 87.590 220.720 89.970 221.525 ;
        RECT 90.810 220.720 93.190 221.525 ;
        RECT 94.030 220.720 102.850 221.525 ;
        RECT 103.690 220.720 112.510 221.525 ;
        RECT 113.350 220.720 115.730 221.525 ;
        RECT 116.570 220.720 118.950 221.525 ;
        RECT 119.790 220.720 131.830 221.525 ;
        RECT 132.670 220.720 160.810 221.525 ;
        RECT 161.650 220.720 199.450 221.525 ;
        RECT 200.290 220.720 202.670 221.525 ;
        RECT 203.510 220.720 205.890 221.525 ;
        RECT 206.730 220.720 217.950 221.525 ;
        RECT 4.230 4.280 217.950 220.720 ;
        RECT 4.230 4.000 70.650 4.280 ;
        RECT 71.490 4.000 80.310 4.280 ;
        RECT 81.150 4.000 83.530 4.280 ;
        RECT 84.370 4.000 86.750 4.280 ;
        RECT 87.590 4.000 89.970 4.280 ;
        RECT 90.810 4.000 93.190 4.280 ;
        RECT 94.030 4.000 109.290 4.280 ;
        RECT 110.130 4.000 217.950 4.280 ;
      LAYER met3 ;
        RECT 3.990 205.040 221.000 221.505 ;
        RECT 3.990 203.640 220.600 205.040 ;
        RECT 3.990 198.240 221.000 203.640 ;
        RECT 3.990 196.840 220.600 198.240 ;
        RECT 3.990 191.440 221.000 196.840 ;
        RECT 4.400 190.040 221.000 191.440 ;
        RECT 3.990 188.040 221.000 190.040 ;
        RECT 4.400 186.640 220.600 188.040 ;
        RECT 3.990 174.440 221.000 186.640 ;
        RECT 3.990 173.040 220.600 174.440 ;
        RECT 3.990 160.840 221.000 173.040 ;
        RECT 3.990 159.440 220.600 160.840 ;
        RECT 3.990 154.040 221.000 159.440 ;
        RECT 4.400 152.640 220.600 154.040 ;
        RECT 3.990 150.640 221.000 152.640 ;
        RECT 3.990 149.240 220.600 150.640 ;
        RECT 3.990 143.840 221.000 149.240 ;
        RECT 3.990 142.440 220.600 143.840 ;
        RECT 3.990 140.440 221.000 142.440 ;
        RECT 4.400 139.040 220.600 140.440 ;
        RECT 3.990 137.040 221.000 139.040 ;
        RECT 3.990 135.640 220.600 137.040 ;
        RECT 3.990 130.240 221.000 135.640 ;
        RECT 3.990 128.840 220.600 130.240 ;
        RECT 3.990 126.840 221.000 128.840 ;
        RECT 3.990 125.440 220.600 126.840 ;
        RECT 3.990 123.440 221.000 125.440 ;
        RECT 4.400 122.040 221.000 123.440 ;
        RECT 3.990 120.040 221.000 122.040 ;
        RECT 4.400 118.640 220.600 120.040 ;
        RECT 3.990 116.640 221.000 118.640 ;
        RECT 4.400 115.240 221.000 116.640 ;
        RECT 3.990 113.240 221.000 115.240 ;
        RECT 4.400 111.840 221.000 113.240 ;
        RECT 3.990 109.840 221.000 111.840 ;
        RECT 4.400 108.440 221.000 109.840 ;
        RECT 3.990 106.440 221.000 108.440 ;
        RECT 4.400 105.040 221.000 106.440 ;
        RECT 3.990 103.040 221.000 105.040 ;
        RECT 4.400 101.640 221.000 103.040 ;
        RECT 3.990 99.640 221.000 101.640 ;
        RECT 4.400 98.240 221.000 99.640 ;
        RECT 3.990 96.240 221.000 98.240 ;
        RECT 4.400 94.840 221.000 96.240 ;
        RECT 3.990 92.840 221.000 94.840 ;
        RECT 4.400 91.440 221.000 92.840 ;
        RECT 3.990 89.440 221.000 91.440 ;
        RECT 4.400 88.040 221.000 89.440 ;
        RECT 3.990 86.040 221.000 88.040 ;
        RECT 4.400 84.640 221.000 86.040 ;
        RECT 3.990 82.640 221.000 84.640 ;
        RECT 4.400 81.240 221.000 82.640 ;
        RECT 3.990 79.240 221.000 81.240 ;
        RECT 4.400 77.840 221.000 79.240 ;
        RECT 3.990 75.840 221.000 77.840 ;
        RECT 4.400 74.440 221.000 75.840 ;
        RECT 3.990 72.440 221.000 74.440 ;
        RECT 4.400 71.040 221.000 72.440 ;
        RECT 3.990 69.040 221.000 71.040 ;
        RECT 4.400 67.640 221.000 69.040 ;
        RECT 3.990 65.640 221.000 67.640 ;
        RECT 4.400 64.240 221.000 65.640 ;
        RECT 3.990 62.240 221.000 64.240 ;
        RECT 4.400 60.840 221.000 62.240 ;
        RECT 3.990 58.840 221.000 60.840 ;
        RECT 4.400 57.440 221.000 58.840 ;
        RECT 3.990 10.715 221.000 57.440 ;
      LAYER met4 ;
        RECT 19.615 212.800 191.985 221.505 ;
        RECT 19.615 23.295 20.640 212.800 ;
        RECT 23.040 23.295 23.940 212.800 ;
        RECT 26.340 23.295 174.240 212.800 ;
        RECT 176.640 23.295 177.540 212.800 ;
        RECT 179.940 23.295 191.985 212.800 ;
  END
END mult_16x16
END LIBRARY

