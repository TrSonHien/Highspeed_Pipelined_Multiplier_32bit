VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 415.845 BY 426.565 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 10.640 75.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 10.640 125.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 10.640 175.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 10.640 225.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 10.640 275.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 410.560 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.030 410.560 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 130.030 410.560 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 180.030 410.560 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 230.030 410.560 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 280.030 410.560 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 330.030 410.560 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 410.560 381.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 410.560 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 410.560 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 126.730 410.560 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 176.730 410.560 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 226.730 410.560 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 276.730 410.560 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.730 410.560 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 410.560 378.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 40.840 415.845 41.440 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 95.240 415.845 95.840 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 100.680 415.845 101.280 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 106.120 415.845 106.720 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 111.560 415.845 112.160 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 117.000 415.845 117.600 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 122.440 415.845 123.040 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 127.880 415.845 128.480 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 133.320 415.845 133.920 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 138.760 415.845 139.360 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 144.200 415.845 144.800 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 46.280 415.845 46.880 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 149.640 415.845 150.240 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 155.080 415.845 155.680 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 160.520 415.845 161.120 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 165.960 415.845 166.560 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 171.400 415.845 172.000 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 176.840 415.845 177.440 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 182.280 415.845 182.880 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 187.720 415.845 188.320 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 193.160 415.845 193.760 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 198.600 415.845 199.200 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 51.720 415.845 52.320 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 204.040 415.845 204.640 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 209.480 415.845 210.080 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 214.920 415.845 215.520 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 220.360 415.845 220.960 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 225.800 415.845 226.400 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 231.240 415.845 231.840 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 236.680 415.845 237.280 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 242.120 415.845 242.720 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 247.560 415.845 248.160 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 253.000 415.845 253.600 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 57.160 415.845 57.760 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 258.440 415.845 259.040 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 263.880 415.845 264.480 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 269.320 415.845 269.920 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 274.760 415.845 275.360 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 280.200 415.845 280.800 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 285.640 415.845 286.240 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 291.080 415.845 291.680 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 296.520 415.845 297.120 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 301.960 415.845 302.560 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 307.400 415.845 308.000 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 62.600 415.845 63.200 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 312.840 415.845 313.440 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 318.280 415.845 318.880 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 323.720 415.845 324.320 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 329.160 415.845 329.760 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 334.600 415.845 335.200 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 340.040 415.845 340.640 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 345.480 415.845 346.080 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 350.920 415.845 351.520 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 356.360 415.845 356.960 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 361.800 415.845 362.400 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 68.040 415.845 68.640 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 367.240 415.845 367.840 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 372.680 415.845 373.280 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 378.120 415.845 378.720 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 383.560 415.845 384.160 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 73.480 415.845 74.080 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 78.920 415.845 79.520 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 84.360 415.845 84.960 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 89.800 415.845 90.400 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 410.510 413.525 ;
      LAYER li1 ;
        RECT 5.520 10.795 410.320 413.525 ;
      LAYER met1 ;
        RECT 3.750 6.840 410.620 414.080 ;
      LAYER met2 ;
        RECT 3.770 4.280 410.220 414.110 ;
        RECT 3.770 0.155 8.550 4.280 ;
        RECT 9.390 0.155 20.970 4.280 ;
        RECT 21.810 0.155 33.390 4.280 ;
        RECT 34.230 0.155 45.810 4.280 ;
        RECT 46.650 0.155 58.230 4.280 ;
        RECT 59.070 0.155 70.650 4.280 ;
        RECT 71.490 0.155 83.070 4.280 ;
        RECT 83.910 0.155 95.490 4.280 ;
        RECT 96.330 0.155 107.910 4.280 ;
        RECT 108.750 0.155 120.330 4.280 ;
        RECT 121.170 0.155 132.750 4.280 ;
        RECT 133.590 0.155 145.170 4.280 ;
        RECT 146.010 0.155 157.590 4.280 ;
        RECT 158.430 0.155 170.010 4.280 ;
        RECT 170.850 0.155 182.430 4.280 ;
        RECT 183.270 0.155 194.850 4.280 ;
        RECT 195.690 0.155 207.270 4.280 ;
        RECT 208.110 0.155 219.690 4.280 ;
        RECT 220.530 0.155 232.110 4.280 ;
        RECT 232.950 0.155 244.530 4.280 ;
        RECT 245.370 0.155 256.950 4.280 ;
        RECT 257.790 0.155 269.370 4.280 ;
        RECT 270.210 0.155 281.790 4.280 ;
        RECT 282.630 0.155 294.210 4.280 ;
        RECT 295.050 0.155 306.630 4.280 ;
        RECT 307.470 0.155 319.050 4.280 ;
        RECT 319.890 0.155 331.470 4.280 ;
        RECT 332.310 0.155 343.890 4.280 ;
        RECT 344.730 0.155 356.310 4.280 ;
        RECT 357.150 0.155 368.730 4.280 ;
        RECT 369.570 0.155 381.150 4.280 ;
        RECT 381.990 0.155 393.570 4.280 ;
        RECT 394.410 0.155 405.990 4.280 ;
        RECT 406.830 0.155 410.220 4.280 ;
      LAYER met3 ;
        RECT 3.745 409.040 411.845 413.605 ;
        RECT 4.400 407.640 411.845 409.040 ;
        RECT 3.745 396.800 411.845 407.640 ;
        RECT 4.400 395.400 411.845 396.800 ;
        RECT 3.745 384.560 411.845 395.400 ;
        RECT 4.400 383.160 411.445 384.560 ;
        RECT 3.745 379.120 411.845 383.160 ;
        RECT 3.745 377.720 411.445 379.120 ;
        RECT 3.745 373.680 411.845 377.720 ;
        RECT 3.745 372.320 411.445 373.680 ;
        RECT 4.400 372.280 411.445 372.320 ;
        RECT 4.400 370.920 411.845 372.280 ;
        RECT 3.745 368.240 411.845 370.920 ;
        RECT 3.745 366.840 411.445 368.240 ;
        RECT 3.745 362.800 411.845 366.840 ;
        RECT 3.745 361.400 411.445 362.800 ;
        RECT 3.745 360.080 411.845 361.400 ;
        RECT 4.400 358.680 411.845 360.080 ;
        RECT 3.745 357.360 411.845 358.680 ;
        RECT 3.745 355.960 411.445 357.360 ;
        RECT 3.745 351.920 411.845 355.960 ;
        RECT 3.745 350.520 411.445 351.920 ;
        RECT 3.745 347.840 411.845 350.520 ;
        RECT 4.400 346.480 411.845 347.840 ;
        RECT 4.400 346.440 411.445 346.480 ;
        RECT 3.745 345.080 411.445 346.440 ;
        RECT 3.745 341.040 411.845 345.080 ;
        RECT 3.745 339.640 411.445 341.040 ;
        RECT 3.745 335.600 411.845 339.640 ;
        RECT 4.400 334.200 411.445 335.600 ;
        RECT 3.745 330.160 411.845 334.200 ;
        RECT 3.745 328.760 411.445 330.160 ;
        RECT 3.745 324.720 411.845 328.760 ;
        RECT 3.745 323.360 411.445 324.720 ;
        RECT 4.400 323.320 411.445 323.360 ;
        RECT 4.400 321.960 411.845 323.320 ;
        RECT 3.745 319.280 411.845 321.960 ;
        RECT 3.745 317.880 411.445 319.280 ;
        RECT 3.745 313.840 411.845 317.880 ;
        RECT 3.745 312.440 411.445 313.840 ;
        RECT 3.745 311.120 411.845 312.440 ;
        RECT 4.400 309.720 411.845 311.120 ;
        RECT 3.745 308.400 411.845 309.720 ;
        RECT 3.745 307.000 411.445 308.400 ;
        RECT 3.745 302.960 411.845 307.000 ;
        RECT 3.745 301.560 411.445 302.960 ;
        RECT 3.745 298.880 411.845 301.560 ;
        RECT 4.400 297.520 411.845 298.880 ;
        RECT 4.400 297.480 411.445 297.520 ;
        RECT 3.745 296.120 411.445 297.480 ;
        RECT 3.745 292.080 411.845 296.120 ;
        RECT 3.745 290.680 411.445 292.080 ;
        RECT 3.745 286.640 411.845 290.680 ;
        RECT 4.400 285.240 411.445 286.640 ;
        RECT 3.745 281.200 411.845 285.240 ;
        RECT 3.745 279.800 411.445 281.200 ;
        RECT 3.745 275.760 411.845 279.800 ;
        RECT 3.745 274.400 411.445 275.760 ;
        RECT 4.400 274.360 411.445 274.400 ;
        RECT 4.400 273.000 411.845 274.360 ;
        RECT 3.745 270.320 411.845 273.000 ;
        RECT 3.745 268.920 411.445 270.320 ;
        RECT 3.745 264.880 411.845 268.920 ;
        RECT 3.745 263.480 411.445 264.880 ;
        RECT 3.745 262.160 411.845 263.480 ;
        RECT 4.400 260.760 411.845 262.160 ;
        RECT 3.745 259.440 411.845 260.760 ;
        RECT 3.745 258.040 411.445 259.440 ;
        RECT 3.745 254.000 411.845 258.040 ;
        RECT 3.745 252.600 411.445 254.000 ;
        RECT 3.745 249.920 411.845 252.600 ;
        RECT 4.400 248.560 411.845 249.920 ;
        RECT 4.400 248.520 411.445 248.560 ;
        RECT 3.745 247.160 411.445 248.520 ;
        RECT 3.745 243.120 411.845 247.160 ;
        RECT 3.745 241.720 411.445 243.120 ;
        RECT 3.745 237.680 411.845 241.720 ;
        RECT 4.400 236.280 411.445 237.680 ;
        RECT 3.745 232.240 411.845 236.280 ;
        RECT 3.745 230.840 411.445 232.240 ;
        RECT 3.745 226.800 411.845 230.840 ;
        RECT 3.745 225.440 411.445 226.800 ;
        RECT 4.400 225.400 411.445 225.440 ;
        RECT 4.400 224.040 411.845 225.400 ;
        RECT 3.745 221.360 411.845 224.040 ;
        RECT 3.745 219.960 411.445 221.360 ;
        RECT 3.745 215.920 411.845 219.960 ;
        RECT 3.745 214.520 411.445 215.920 ;
        RECT 3.745 213.200 411.845 214.520 ;
        RECT 4.400 211.800 411.845 213.200 ;
        RECT 3.745 210.480 411.845 211.800 ;
        RECT 3.745 209.080 411.445 210.480 ;
        RECT 3.745 205.040 411.845 209.080 ;
        RECT 3.745 203.640 411.445 205.040 ;
        RECT 3.745 200.960 411.845 203.640 ;
        RECT 4.400 199.600 411.845 200.960 ;
        RECT 4.400 199.560 411.445 199.600 ;
        RECT 3.745 198.200 411.445 199.560 ;
        RECT 3.745 194.160 411.845 198.200 ;
        RECT 3.745 192.760 411.445 194.160 ;
        RECT 3.745 188.720 411.845 192.760 ;
        RECT 4.400 187.320 411.445 188.720 ;
        RECT 3.745 183.280 411.845 187.320 ;
        RECT 3.745 181.880 411.445 183.280 ;
        RECT 3.745 177.840 411.845 181.880 ;
        RECT 3.745 176.480 411.445 177.840 ;
        RECT 4.400 176.440 411.445 176.480 ;
        RECT 4.400 175.080 411.845 176.440 ;
        RECT 3.745 172.400 411.845 175.080 ;
        RECT 3.745 171.000 411.445 172.400 ;
        RECT 3.745 166.960 411.845 171.000 ;
        RECT 3.745 165.560 411.445 166.960 ;
        RECT 3.745 164.240 411.845 165.560 ;
        RECT 4.400 162.840 411.845 164.240 ;
        RECT 3.745 161.520 411.845 162.840 ;
        RECT 3.745 160.120 411.445 161.520 ;
        RECT 3.745 156.080 411.845 160.120 ;
        RECT 3.745 154.680 411.445 156.080 ;
        RECT 3.745 152.000 411.845 154.680 ;
        RECT 4.400 150.640 411.845 152.000 ;
        RECT 4.400 150.600 411.445 150.640 ;
        RECT 3.745 149.240 411.445 150.600 ;
        RECT 3.745 145.200 411.845 149.240 ;
        RECT 3.745 143.800 411.445 145.200 ;
        RECT 3.745 139.760 411.845 143.800 ;
        RECT 4.400 138.360 411.445 139.760 ;
        RECT 3.745 134.320 411.845 138.360 ;
        RECT 3.745 132.920 411.445 134.320 ;
        RECT 3.745 128.880 411.845 132.920 ;
        RECT 3.745 127.520 411.445 128.880 ;
        RECT 4.400 127.480 411.445 127.520 ;
        RECT 4.400 126.120 411.845 127.480 ;
        RECT 3.745 123.440 411.845 126.120 ;
        RECT 3.745 122.040 411.445 123.440 ;
        RECT 3.745 118.000 411.845 122.040 ;
        RECT 3.745 116.600 411.445 118.000 ;
        RECT 3.745 115.280 411.845 116.600 ;
        RECT 4.400 113.880 411.845 115.280 ;
        RECT 3.745 112.560 411.845 113.880 ;
        RECT 3.745 111.160 411.445 112.560 ;
        RECT 3.745 107.120 411.845 111.160 ;
        RECT 3.745 105.720 411.445 107.120 ;
        RECT 3.745 103.040 411.845 105.720 ;
        RECT 4.400 101.680 411.845 103.040 ;
        RECT 4.400 101.640 411.445 101.680 ;
        RECT 3.745 100.280 411.445 101.640 ;
        RECT 3.745 96.240 411.845 100.280 ;
        RECT 3.745 94.840 411.445 96.240 ;
        RECT 3.745 90.800 411.845 94.840 ;
        RECT 4.400 89.400 411.445 90.800 ;
        RECT 3.745 85.360 411.845 89.400 ;
        RECT 3.745 83.960 411.445 85.360 ;
        RECT 3.745 79.920 411.845 83.960 ;
        RECT 3.745 78.560 411.445 79.920 ;
        RECT 4.400 78.520 411.445 78.560 ;
        RECT 4.400 77.160 411.845 78.520 ;
        RECT 3.745 74.480 411.845 77.160 ;
        RECT 3.745 73.080 411.445 74.480 ;
        RECT 3.745 69.040 411.845 73.080 ;
        RECT 3.745 67.640 411.445 69.040 ;
        RECT 3.745 66.320 411.845 67.640 ;
        RECT 4.400 64.920 411.845 66.320 ;
        RECT 3.745 63.600 411.845 64.920 ;
        RECT 3.745 62.200 411.445 63.600 ;
        RECT 3.745 58.160 411.845 62.200 ;
        RECT 3.745 56.760 411.445 58.160 ;
        RECT 3.745 54.080 411.845 56.760 ;
        RECT 4.400 52.720 411.845 54.080 ;
        RECT 4.400 52.680 411.445 52.720 ;
        RECT 3.745 51.320 411.445 52.680 ;
        RECT 3.745 47.280 411.845 51.320 ;
        RECT 3.745 45.880 411.445 47.280 ;
        RECT 3.745 41.840 411.845 45.880 ;
        RECT 4.400 40.440 411.445 41.840 ;
        RECT 3.745 29.600 411.845 40.440 ;
        RECT 4.400 28.200 411.845 29.600 ;
        RECT 3.745 17.360 411.845 28.200 ;
        RECT 4.400 15.960 411.845 17.360 ;
        RECT 3.745 0.175 411.845 15.960 ;
      LAYER met4 ;
        RECT 3.975 10.240 20.640 402.385 ;
        RECT 23.040 10.240 23.940 402.385 ;
        RECT 26.340 10.240 70.640 402.385 ;
        RECT 73.040 10.240 73.940 402.385 ;
        RECT 76.340 10.240 120.640 402.385 ;
        RECT 123.040 10.240 123.940 402.385 ;
        RECT 126.340 10.240 170.640 402.385 ;
        RECT 173.040 10.240 173.940 402.385 ;
        RECT 176.340 10.240 220.640 402.385 ;
        RECT 223.040 10.240 223.940 402.385 ;
        RECT 226.340 10.240 270.640 402.385 ;
        RECT 273.040 10.240 273.940 402.385 ;
        RECT 276.340 10.240 320.640 402.385 ;
        RECT 323.040 10.240 323.940 402.385 ;
        RECT 326.340 10.240 370.640 402.385 ;
        RECT 373.040 10.240 373.940 402.385 ;
        RECT 376.340 10.240 390.705 402.385 ;
        RECT 3.975 0.175 390.705 10.240 ;
  END
END pipelined_mult
END LIBRARY

