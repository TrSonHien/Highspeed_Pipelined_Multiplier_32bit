VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 10.640 75.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 10.640 125.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 10.640 175.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 10.640 225.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 10.640 275.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.340 10.640 475.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.340 10.640 525.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.340 10.640 575.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 624.340 10.640 625.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 674.340 10.640 675.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 724.340 10.640 725.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 774.340 10.640 775.940 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 794.660 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.030 794.660 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 130.030 794.660 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 180.030 794.660 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 230.030 794.660 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 280.030 794.660 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 330.030 794.660 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 794.660 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 430.030 794.660 431.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 480.030 794.660 481.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 530.030 794.660 531.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 580.030 794.660 581.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 630.030 794.660 631.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 680.030 794.660 681.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 730.030 794.660 731.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 780.030 794.660 781.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 789.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 794.660 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 794.660 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 126.730 794.660 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 176.730 794.660 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 226.730 794.660 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 276.730 794.660 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.730 794.660 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 794.660 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 426.730 794.660 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 476.730 794.660 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 526.730 794.660 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 576.730 794.660 578.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 626.730 794.660 628.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 676.730 794.660 678.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 726.730 794.660 728.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 776.730 794.660 778.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 745.320 4.000 745.920 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 543.350 0.000 543.630 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 662.950 0.000 663.230 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 734.710 0.000 734.990 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 557.640 800.000 558.240 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 312.840 800.000 313.440 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 337.320 800.000 337.920 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 361.800 800.000 362.400 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 386.280 800.000 386.880 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 410.760 800.000 411.360 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 435.240 800.000 435.840 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.720 800.000 460.320 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 484.200 800.000 484.800 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 508.680 800.000 509.280 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 533.160 800.000 533.760 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 582.120 800.000 582.720 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 68.040 800.000 68.640 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 92.520 800.000 93.120 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 117.000 800.000 117.600 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 141.480 800.000 142.080 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 165.960 800.000 166.560 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 190.440 800.000 191.040 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 214.920 800.000 215.520 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 239.400 800.000 240.000 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 263.880 800.000 264.480 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 288.360 800.000 288.960 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 606.600 800.000 607.200 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 19.080 800.000 19.680 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 43.560 800.000 44.160 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 610.970 796.000 611.250 800.000 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 635.810 796.000 636.090 800.000 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 660.650 796.000 660.930 800.000 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 685.490 796.000 685.770 800.000 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 710.330 796.000 710.610 800.000 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 735.170 796.000 735.450 800.000 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 760.010 796.000 760.290 800.000 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 784.850 796.000 785.130 800.000 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 631.080 800.000 631.680 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 362.570 796.000 362.850 800.000 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 387.410 796.000 387.690 800.000 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 796.000 412.530 800.000 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 437.090 796.000 437.370 800.000 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 461.930 796.000 462.210 800.000 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 486.770 796.000 487.050 800.000 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 511.610 796.000 511.890 800.000 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 536.450 796.000 536.730 800.000 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 561.290 796.000 561.570 800.000 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 586.130 796.000 586.410 800.000 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 655.560 800.000 656.160 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 796.000 114.450 800.000 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.010 796.000 139.290 800.000 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 163.850 796.000 164.130 800.000 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.690 796.000 188.970 800.000 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 213.530 796.000 213.810 800.000 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 796.000 238.650 800.000 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 263.210 796.000 263.490 800.000 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 288.050 796.000 288.330 800.000 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 312.890 796.000 313.170 800.000 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 337.730 796.000 338.010 800.000 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 680.040 800.000 680.640 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 14.810 796.000 15.090 800.000 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 796.000 39.930 800.000 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 796.000 64.770 800.000 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 89.330 796.000 89.610 800.000 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 704.520 800.000 705.120 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 729.000 800.000 729.600 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 753.480 800.000 754.080 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 777.960 800.000 778.560 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 794.610 788.885 ;
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 4.210 10.640 794.420 789.040 ;
      LAYER met2 ;
        RECT 4.230 795.720 14.530 796.690 ;
        RECT 15.370 795.720 39.370 796.690 ;
        RECT 40.210 795.720 64.210 796.690 ;
        RECT 65.050 795.720 89.050 796.690 ;
        RECT 89.890 795.720 113.890 796.690 ;
        RECT 114.730 795.720 138.730 796.690 ;
        RECT 139.570 795.720 163.570 796.690 ;
        RECT 164.410 795.720 188.410 796.690 ;
        RECT 189.250 795.720 213.250 796.690 ;
        RECT 214.090 795.720 238.090 796.690 ;
        RECT 238.930 795.720 262.930 796.690 ;
        RECT 263.770 795.720 287.770 796.690 ;
        RECT 288.610 795.720 312.610 796.690 ;
        RECT 313.450 795.720 337.450 796.690 ;
        RECT 338.290 795.720 362.290 796.690 ;
        RECT 363.130 795.720 387.130 796.690 ;
        RECT 387.970 795.720 411.970 796.690 ;
        RECT 412.810 795.720 436.810 796.690 ;
        RECT 437.650 795.720 461.650 796.690 ;
        RECT 462.490 795.720 486.490 796.690 ;
        RECT 487.330 795.720 511.330 796.690 ;
        RECT 512.170 795.720 536.170 796.690 ;
        RECT 537.010 795.720 561.010 796.690 ;
        RECT 561.850 795.720 585.850 796.690 ;
        RECT 586.690 795.720 610.690 796.690 ;
        RECT 611.530 795.720 635.530 796.690 ;
        RECT 636.370 795.720 660.370 796.690 ;
        RECT 661.210 795.720 685.210 796.690 ;
        RECT 686.050 795.720 710.050 796.690 ;
        RECT 710.890 795.720 734.890 796.690 ;
        RECT 735.730 795.720 759.730 796.690 ;
        RECT 760.570 795.720 784.570 796.690 ;
        RECT 785.410 795.720 792.940 796.690 ;
        RECT 4.230 4.280 792.940 795.720 ;
        RECT 4.230 4.000 16.830 4.280 ;
        RECT 17.670 4.000 40.750 4.280 ;
        RECT 41.590 4.000 64.670 4.280 ;
        RECT 65.510 4.000 88.590 4.280 ;
        RECT 89.430 4.000 112.510 4.280 ;
        RECT 113.350 4.000 136.430 4.280 ;
        RECT 137.270 4.000 160.350 4.280 ;
        RECT 161.190 4.000 184.270 4.280 ;
        RECT 185.110 4.000 208.190 4.280 ;
        RECT 209.030 4.000 232.110 4.280 ;
        RECT 232.950 4.000 256.030 4.280 ;
        RECT 256.870 4.000 279.950 4.280 ;
        RECT 280.790 4.000 303.870 4.280 ;
        RECT 304.710 4.000 327.790 4.280 ;
        RECT 328.630 4.000 351.710 4.280 ;
        RECT 352.550 4.000 375.630 4.280 ;
        RECT 376.470 4.000 399.550 4.280 ;
        RECT 400.390 4.000 423.470 4.280 ;
        RECT 424.310 4.000 447.390 4.280 ;
        RECT 448.230 4.000 471.310 4.280 ;
        RECT 472.150 4.000 495.230 4.280 ;
        RECT 496.070 4.000 519.150 4.280 ;
        RECT 519.990 4.000 543.070 4.280 ;
        RECT 543.910 4.000 566.990 4.280 ;
        RECT 567.830 4.000 590.910 4.280 ;
        RECT 591.750 4.000 614.830 4.280 ;
        RECT 615.670 4.000 638.750 4.280 ;
        RECT 639.590 4.000 662.670 4.280 ;
        RECT 663.510 4.000 686.590 4.280 ;
        RECT 687.430 4.000 710.510 4.280 ;
        RECT 711.350 4.000 734.430 4.280 ;
        RECT 735.270 4.000 758.350 4.280 ;
        RECT 759.190 4.000 782.270 4.280 ;
        RECT 783.110 4.000 792.940 4.280 ;
      LAYER met3 ;
        RECT 3.990 778.960 796.000 788.965 ;
        RECT 3.990 777.560 795.600 778.960 ;
        RECT 3.990 769.440 796.000 777.560 ;
        RECT 4.400 768.040 796.000 769.440 ;
        RECT 3.990 754.480 796.000 768.040 ;
        RECT 3.990 753.080 795.600 754.480 ;
        RECT 3.990 746.320 796.000 753.080 ;
        RECT 4.400 744.920 796.000 746.320 ;
        RECT 3.990 730.000 796.000 744.920 ;
        RECT 3.990 728.600 795.600 730.000 ;
        RECT 3.990 723.200 796.000 728.600 ;
        RECT 4.400 721.800 796.000 723.200 ;
        RECT 3.990 705.520 796.000 721.800 ;
        RECT 3.990 704.120 795.600 705.520 ;
        RECT 3.990 700.080 796.000 704.120 ;
        RECT 4.400 698.680 796.000 700.080 ;
        RECT 3.990 681.040 796.000 698.680 ;
        RECT 3.990 679.640 795.600 681.040 ;
        RECT 3.990 676.960 796.000 679.640 ;
        RECT 4.400 675.560 796.000 676.960 ;
        RECT 3.990 656.560 796.000 675.560 ;
        RECT 3.990 655.160 795.600 656.560 ;
        RECT 3.990 653.840 796.000 655.160 ;
        RECT 4.400 652.440 796.000 653.840 ;
        RECT 3.990 632.080 796.000 652.440 ;
        RECT 3.990 630.720 795.600 632.080 ;
        RECT 4.400 630.680 795.600 630.720 ;
        RECT 4.400 629.320 796.000 630.680 ;
        RECT 3.990 607.600 796.000 629.320 ;
        RECT 4.400 606.200 795.600 607.600 ;
        RECT 3.990 584.480 796.000 606.200 ;
        RECT 4.400 583.120 796.000 584.480 ;
        RECT 4.400 583.080 795.600 583.120 ;
        RECT 3.990 581.720 795.600 583.080 ;
        RECT 3.990 561.360 796.000 581.720 ;
        RECT 4.400 559.960 796.000 561.360 ;
        RECT 3.990 558.640 796.000 559.960 ;
        RECT 3.990 557.240 795.600 558.640 ;
        RECT 3.990 538.240 796.000 557.240 ;
        RECT 4.400 536.840 796.000 538.240 ;
        RECT 3.990 534.160 796.000 536.840 ;
        RECT 3.990 532.760 795.600 534.160 ;
        RECT 3.990 515.120 796.000 532.760 ;
        RECT 4.400 513.720 796.000 515.120 ;
        RECT 3.990 509.680 796.000 513.720 ;
        RECT 3.990 508.280 795.600 509.680 ;
        RECT 3.990 492.000 796.000 508.280 ;
        RECT 4.400 490.600 796.000 492.000 ;
        RECT 3.990 485.200 796.000 490.600 ;
        RECT 3.990 483.800 795.600 485.200 ;
        RECT 3.990 468.880 796.000 483.800 ;
        RECT 4.400 467.480 796.000 468.880 ;
        RECT 3.990 460.720 796.000 467.480 ;
        RECT 3.990 459.320 795.600 460.720 ;
        RECT 3.990 445.760 796.000 459.320 ;
        RECT 4.400 444.360 796.000 445.760 ;
        RECT 3.990 436.240 796.000 444.360 ;
        RECT 3.990 434.840 795.600 436.240 ;
        RECT 3.990 422.640 796.000 434.840 ;
        RECT 4.400 421.240 796.000 422.640 ;
        RECT 3.990 411.760 796.000 421.240 ;
        RECT 3.990 410.360 795.600 411.760 ;
        RECT 3.990 399.520 796.000 410.360 ;
        RECT 4.400 398.120 796.000 399.520 ;
        RECT 3.990 387.280 796.000 398.120 ;
        RECT 3.990 385.880 795.600 387.280 ;
        RECT 3.990 376.400 796.000 385.880 ;
        RECT 4.400 375.000 796.000 376.400 ;
        RECT 3.990 362.800 796.000 375.000 ;
        RECT 3.990 361.400 795.600 362.800 ;
        RECT 3.990 353.280 796.000 361.400 ;
        RECT 4.400 351.880 796.000 353.280 ;
        RECT 3.990 338.320 796.000 351.880 ;
        RECT 3.990 336.920 795.600 338.320 ;
        RECT 3.990 330.160 796.000 336.920 ;
        RECT 4.400 328.760 796.000 330.160 ;
        RECT 3.990 313.840 796.000 328.760 ;
        RECT 3.990 312.440 795.600 313.840 ;
        RECT 3.990 307.040 796.000 312.440 ;
        RECT 4.400 305.640 796.000 307.040 ;
        RECT 3.990 289.360 796.000 305.640 ;
        RECT 3.990 287.960 795.600 289.360 ;
        RECT 3.990 283.920 796.000 287.960 ;
        RECT 4.400 282.520 796.000 283.920 ;
        RECT 3.990 264.880 796.000 282.520 ;
        RECT 3.990 263.480 795.600 264.880 ;
        RECT 3.990 260.800 796.000 263.480 ;
        RECT 4.400 259.400 796.000 260.800 ;
        RECT 3.990 240.400 796.000 259.400 ;
        RECT 3.990 239.000 795.600 240.400 ;
        RECT 3.990 237.680 796.000 239.000 ;
        RECT 4.400 236.280 796.000 237.680 ;
        RECT 3.990 215.920 796.000 236.280 ;
        RECT 3.990 214.560 795.600 215.920 ;
        RECT 4.400 214.520 795.600 214.560 ;
        RECT 4.400 213.160 796.000 214.520 ;
        RECT 3.990 191.440 796.000 213.160 ;
        RECT 4.400 190.040 795.600 191.440 ;
        RECT 3.990 168.320 796.000 190.040 ;
        RECT 4.400 166.960 796.000 168.320 ;
        RECT 4.400 166.920 795.600 166.960 ;
        RECT 3.990 165.560 795.600 166.920 ;
        RECT 3.990 145.200 796.000 165.560 ;
        RECT 4.400 143.800 796.000 145.200 ;
        RECT 3.990 142.480 796.000 143.800 ;
        RECT 3.990 141.080 795.600 142.480 ;
        RECT 3.990 122.080 796.000 141.080 ;
        RECT 4.400 120.680 796.000 122.080 ;
        RECT 3.990 118.000 796.000 120.680 ;
        RECT 3.990 116.600 795.600 118.000 ;
        RECT 3.990 98.960 796.000 116.600 ;
        RECT 4.400 97.560 796.000 98.960 ;
        RECT 3.990 93.520 796.000 97.560 ;
        RECT 3.990 92.120 795.600 93.520 ;
        RECT 3.990 75.840 796.000 92.120 ;
        RECT 4.400 74.440 796.000 75.840 ;
        RECT 3.990 69.040 796.000 74.440 ;
        RECT 3.990 67.640 795.600 69.040 ;
        RECT 3.990 52.720 796.000 67.640 ;
        RECT 4.400 51.320 796.000 52.720 ;
        RECT 3.990 44.560 796.000 51.320 ;
        RECT 3.990 43.160 795.600 44.560 ;
        RECT 3.990 29.600 796.000 43.160 ;
        RECT 4.400 28.200 796.000 29.600 ;
        RECT 3.990 20.080 796.000 28.200 ;
        RECT 3.990 18.680 795.600 20.080 ;
        RECT 3.990 10.715 796.000 18.680 ;
      LAYER met4 ;
        RECT 197.175 13.095 220.640 539.745 ;
        RECT 223.040 13.095 223.940 539.745 ;
        RECT 226.340 13.095 270.640 539.745 ;
        RECT 273.040 13.095 273.940 539.745 ;
        RECT 276.340 13.095 320.640 539.745 ;
        RECT 323.040 13.095 323.940 539.745 ;
        RECT 326.340 13.095 370.640 539.745 ;
        RECT 373.040 13.095 373.940 539.745 ;
        RECT 376.340 13.095 420.640 539.745 ;
        RECT 423.040 13.095 423.940 539.745 ;
        RECT 426.340 13.095 470.640 539.745 ;
        RECT 473.040 13.095 473.940 539.745 ;
        RECT 476.340 13.095 520.640 539.745 ;
        RECT 523.040 13.095 523.940 539.745 ;
        RECT 526.340 13.095 570.640 539.745 ;
        RECT 573.040 13.095 573.940 539.745 ;
        RECT 576.340 13.095 620.640 539.745 ;
        RECT 623.040 13.095 623.940 539.745 ;
        RECT 626.340 13.095 643.705 539.745 ;
      LAYER met5 ;
        RECT 309.700 383.230 591.900 393.500 ;
        RECT 309.700 368.100 591.900 375.130 ;
  END
END pipelined_mult
END LIBRARY

