VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 415.845 BY 426.565 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 10.640 75.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 10.640 125.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 10.640 175.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 10.640 225.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 10.640 275.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 410.560 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.030 410.560 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 130.030 410.560 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 180.030 410.560 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 230.030 410.560 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 280.030 410.560 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 330.030 410.560 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 410.560 381.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 413.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 413.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 410.560 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 410.560 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 126.730 410.560 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 176.730 410.560 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 226.730 410.560 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 276.730 410.560 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.730 410.560 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 410.560 378.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 381.430 0.000 381.710 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 292.440 415.845 293.040 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 170.040 415.845 170.640 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 182.280 415.845 182.880 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 194.520 415.845 195.120 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 206.760 415.845 207.360 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 219.000 415.845 219.600 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 231.240 415.845 231.840 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 243.480 415.845 244.080 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 255.720 415.845 256.320 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 267.960 415.845 268.560 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 280.200 415.845 280.800 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 304.680 415.845 305.280 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 47.640 415.845 48.240 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 59.880 415.845 60.480 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 72.120 415.845 72.720 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 84.360 415.845 84.960 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 96.600 415.845 97.200 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 108.840 415.845 109.440 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 121.080 415.845 121.680 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 133.320 415.845 133.920 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 145.560 415.845 146.160 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 157.800 415.845 158.400 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 316.920 415.845 317.520 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 23.160 415.845 23.760 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 35.400 415.845 36.000 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.030 422.565 317.310 426.565 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 329.910 422.565 330.190 426.565 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 342.790 422.565 343.070 426.565 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 355.670 422.565 355.950 426.565 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 368.550 422.565 368.830 426.565 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 381.430 422.565 381.710 426.565 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 394.310 422.565 394.590 426.565 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 407.190 422.565 407.470 426.565 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 329.160 415.845 329.760 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.230 422.565 188.510 426.565 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 201.110 422.565 201.390 426.565 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 213.990 422.565 214.270 426.565 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 226.870 422.565 227.150 426.565 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 239.750 422.565 240.030 426.565 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 252.630 422.565 252.910 426.565 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 265.510 422.565 265.790 426.565 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 278.390 422.565 278.670 426.565 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 291.270 422.565 291.550 426.565 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 304.150 422.565 304.430 426.565 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 341.400 415.845 342.000 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 422.565 59.710 426.565 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.310 422.565 72.590 426.565 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 85.190 422.565 85.470 426.565 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.070 422.565 98.350 426.565 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.950 422.565 111.230 426.565 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 123.830 422.565 124.110 426.565 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 136.710 422.565 136.990 426.565 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.590 422.565 149.870 426.565 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.470 422.565 162.750 426.565 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.350 422.565 175.630 426.565 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 353.640 415.845 354.240 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 7.910 422.565 8.190 426.565 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 20.790 422.565 21.070 426.565 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 422.565 33.950 426.565 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 422.565 46.830 426.565 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 365.880 415.845 366.480 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 378.120 415.845 378.720 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 390.360 415.845 390.960 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 411.845 402.600 415.845 403.200 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 410.510 413.525 ;
      LAYER li1 ;
        RECT 5.520 10.795 410.320 413.525 ;
      LAYER met1 ;
        RECT 4.210 8.880 410.620 414.080 ;
      LAYER met2 ;
        RECT 4.230 422.285 7.630 423.370 ;
        RECT 8.470 422.285 20.510 423.370 ;
        RECT 21.350 422.285 33.390 423.370 ;
        RECT 34.230 422.285 46.270 423.370 ;
        RECT 47.110 422.285 59.150 423.370 ;
        RECT 59.990 422.285 72.030 423.370 ;
        RECT 72.870 422.285 84.910 423.370 ;
        RECT 85.750 422.285 97.790 423.370 ;
        RECT 98.630 422.285 110.670 423.370 ;
        RECT 111.510 422.285 123.550 423.370 ;
        RECT 124.390 422.285 136.430 423.370 ;
        RECT 137.270 422.285 149.310 423.370 ;
        RECT 150.150 422.285 162.190 423.370 ;
        RECT 163.030 422.285 175.070 423.370 ;
        RECT 175.910 422.285 187.950 423.370 ;
        RECT 188.790 422.285 200.830 423.370 ;
        RECT 201.670 422.285 213.710 423.370 ;
        RECT 214.550 422.285 226.590 423.370 ;
        RECT 227.430 422.285 239.470 423.370 ;
        RECT 240.310 422.285 252.350 423.370 ;
        RECT 253.190 422.285 265.230 423.370 ;
        RECT 266.070 422.285 278.110 423.370 ;
        RECT 278.950 422.285 290.990 423.370 ;
        RECT 291.830 422.285 303.870 423.370 ;
        RECT 304.710 422.285 316.750 423.370 ;
        RECT 317.590 422.285 329.630 423.370 ;
        RECT 330.470 422.285 342.510 423.370 ;
        RECT 343.350 422.285 355.390 423.370 ;
        RECT 356.230 422.285 368.270 423.370 ;
        RECT 369.110 422.285 381.150 423.370 ;
        RECT 381.990 422.285 394.030 423.370 ;
        RECT 394.870 422.285 406.910 423.370 ;
        RECT 407.750 422.285 409.760 423.370 ;
        RECT 4.230 4.280 409.760 422.285 ;
        RECT 4.230 4.000 8.550 4.280 ;
        RECT 9.390 4.000 20.970 4.280 ;
        RECT 21.810 4.000 33.390 4.280 ;
        RECT 34.230 4.000 45.810 4.280 ;
        RECT 46.650 4.000 58.230 4.280 ;
        RECT 59.070 4.000 70.650 4.280 ;
        RECT 71.490 4.000 83.070 4.280 ;
        RECT 83.910 4.000 95.490 4.280 ;
        RECT 96.330 4.000 107.910 4.280 ;
        RECT 108.750 4.000 120.330 4.280 ;
        RECT 121.170 4.000 132.750 4.280 ;
        RECT 133.590 4.000 145.170 4.280 ;
        RECT 146.010 4.000 157.590 4.280 ;
        RECT 158.430 4.000 170.010 4.280 ;
        RECT 170.850 4.000 182.430 4.280 ;
        RECT 183.270 4.000 194.850 4.280 ;
        RECT 195.690 4.000 207.270 4.280 ;
        RECT 208.110 4.000 219.690 4.280 ;
        RECT 220.530 4.000 232.110 4.280 ;
        RECT 232.950 4.000 244.530 4.280 ;
        RECT 245.370 4.000 256.950 4.280 ;
        RECT 257.790 4.000 269.370 4.280 ;
        RECT 270.210 4.000 281.790 4.280 ;
        RECT 282.630 4.000 294.210 4.280 ;
        RECT 295.050 4.000 306.630 4.280 ;
        RECT 307.470 4.000 319.050 4.280 ;
        RECT 319.890 4.000 331.470 4.280 ;
        RECT 332.310 4.000 343.890 4.280 ;
        RECT 344.730 4.000 356.310 4.280 ;
        RECT 357.150 4.000 368.730 4.280 ;
        RECT 369.570 4.000 381.150 4.280 ;
        RECT 381.990 4.000 393.570 4.280 ;
        RECT 394.410 4.000 405.990 4.280 ;
        RECT 406.830 4.000 409.760 4.280 ;
      LAYER met3 ;
        RECT 3.990 409.040 411.845 413.605 ;
        RECT 4.400 407.640 411.845 409.040 ;
        RECT 3.990 403.600 411.845 407.640 ;
        RECT 3.990 402.200 411.445 403.600 ;
        RECT 3.990 396.800 411.845 402.200 ;
        RECT 4.400 395.400 411.845 396.800 ;
        RECT 3.990 391.360 411.845 395.400 ;
        RECT 3.990 389.960 411.445 391.360 ;
        RECT 3.990 384.560 411.845 389.960 ;
        RECT 4.400 383.160 411.845 384.560 ;
        RECT 3.990 379.120 411.845 383.160 ;
        RECT 3.990 377.720 411.445 379.120 ;
        RECT 3.990 372.320 411.845 377.720 ;
        RECT 4.400 370.920 411.845 372.320 ;
        RECT 3.990 366.880 411.845 370.920 ;
        RECT 3.990 365.480 411.445 366.880 ;
        RECT 3.990 360.080 411.845 365.480 ;
        RECT 4.400 358.680 411.845 360.080 ;
        RECT 3.990 354.640 411.845 358.680 ;
        RECT 3.990 353.240 411.445 354.640 ;
        RECT 3.990 347.840 411.845 353.240 ;
        RECT 4.400 346.440 411.845 347.840 ;
        RECT 3.990 342.400 411.845 346.440 ;
        RECT 3.990 341.000 411.445 342.400 ;
        RECT 3.990 335.600 411.845 341.000 ;
        RECT 4.400 334.200 411.845 335.600 ;
        RECT 3.990 330.160 411.845 334.200 ;
        RECT 3.990 328.760 411.445 330.160 ;
        RECT 3.990 323.360 411.845 328.760 ;
        RECT 4.400 321.960 411.845 323.360 ;
        RECT 3.990 317.920 411.845 321.960 ;
        RECT 3.990 316.520 411.445 317.920 ;
        RECT 3.990 311.120 411.845 316.520 ;
        RECT 4.400 309.720 411.845 311.120 ;
        RECT 3.990 305.680 411.845 309.720 ;
        RECT 3.990 304.280 411.445 305.680 ;
        RECT 3.990 298.880 411.845 304.280 ;
        RECT 4.400 297.480 411.845 298.880 ;
        RECT 3.990 293.440 411.845 297.480 ;
        RECT 3.990 292.040 411.445 293.440 ;
        RECT 3.990 286.640 411.845 292.040 ;
        RECT 4.400 285.240 411.845 286.640 ;
        RECT 3.990 281.200 411.845 285.240 ;
        RECT 3.990 279.800 411.445 281.200 ;
        RECT 3.990 274.400 411.845 279.800 ;
        RECT 4.400 273.000 411.845 274.400 ;
        RECT 3.990 268.960 411.845 273.000 ;
        RECT 3.990 267.560 411.445 268.960 ;
        RECT 3.990 262.160 411.845 267.560 ;
        RECT 4.400 260.760 411.845 262.160 ;
        RECT 3.990 256.720 411.845 260.760 ;
        RECT 3.990 255.320 411.445 256.720 ;
        RECT 3.990 249.920 411.845 255.320 ;
        RECT 4.400 248.520 411.845 249.920 ;
        RECT 3.990 244.480 411.845 248.520 ;
        RECT 3.990 243.080 411.445 244.480 ;
        RECT 3.990 237.680 411.845 243.080 ;
        RECT 4.400 236.280 411.845 237.680 ;
        RECT 3.990 232.240 411.845 236.280 ;
        RECT 3.990 230.840 411.445 232.240 ;
        RECT 3.990 225.440 411.845 230.840 ;
        RECT 4.400 224.040 411.845 225.440 ;
        RECT 3.990 220.000 411.845 224.040 ;
        RECT 3.990 218.600 411.445 220.000 ;
        RECT 3.990 213.200 411.845 218.600 ;
        RECT 4.400 211.800 411.845 213.200 ;
        RECT 3.990 207.760 411.845 211.800 ;
        RECT 3.990 206.360 411.445 207.760 ;
        RECT 3.990 200.960 411.845 206.360 ;
        RECT 4.400 199.560 411.845 200.960 ;
        RECT 3.990 195.520 411.845 199.560 ;
        RECT 3.990 194.120 411.445 195.520 ;
        RECT 3.990 188.720 411.845 194.120 ;
        RECT 4.400 187.320 411.845 188.720 ;
        RECT 3.990 183.280 411.845 187.320 ;
        RECT 3.990 181.880 411.445 183.280 ;
        RECT 3.990 176.480 411.845 181.880 ;
        RECT 4.400 175.080 411.845 176.480 ;
        RECT 3.990 171.040 411.845 175.080 ;
        RECT 3.990 169.640 411.445 171.040 ;
        RECT 3.990 164.240 411.845 169.640 ;
        RECT 4.400 162.840 411.845 164.240 ;
        RECT 3.990 158.800 411.845 162.840 ;
        RECT 3.990 157.400 411.445 158.800 ;
        RECT 3.990 152.000 411.845 157.400 ;
        RECT 4.400 150.600 411.845 152.000 ;
        RECT 3.990 146.560 411.845 150.600 ;
        RECT 3.990 145.160 411.445 146.560 ;
        RECT 3.990 139.760 411.845 145.160 ;
        RECT 4.400 138.360 411.845 139.760 ;
        RECT 3.990 134.320 411.845 138.360 ;
        RECT 3.990 132.920 411.445 134.320 ;
        RECT 3.990 127.520 411.845 132.920 ;
        RECT 4.400 126.120 411.845 127.520 ;
        RECT 3.990 122.080 411.845 126.120 ;
        RECT 3.990 120.680 411.445 122.080 ;
        RECT 3.990 115.280 411.845 120.680 ;
        RECT 4.400 113.880 411.845 115.280 ;
        RECT 3.990 109.840 411.845 113.880 ;
        RECT 3.990 108.440 411.445 109.840 ;
        RECT 3.990 103.040 411.845 108.440 ;
        RECT 4.400 101.640 411.845 103.040 ;
        RECT 3.990 97.600 411.845 101.640 ;
        RECT 3.990 96.200 411.445 97.600 ;
        RECT 3.990 90.800 411.845 96.200 ;
        RECT 4.400 89.400 411.845 90.800 ;
        RECT 3.990 85.360 411.845 89.400 ;
        RECT 3.990 83.960 411.445 85.360 ;
        RECT 3.990 78.560 411.845 83.960 ;
        RECT 4.400 77.160 411.845 78.560 ;
        RECT 3.990 73.120 411.845 77.160 ;
        RECT 3.990 71.720 411.445 73.120 ;
        RECT 3.990 66.320 411.845 71.720 ;
        RECT 4.400 64.920 411.845 66.320 ;
        RECT 3.990 60.880 411.845 64.920 ;
        RECT 3.990 59.480 411.445 60.880 ;
        RECT 3.990 54.080 411.845 59.480 ;
        RECT 4.400 52.680 411.845 54.080 ;
        RECT 3.990 48.640 411.845 52.680 ;
        RECT 3.990 47.240 411.445 48.640 ;
        RECT 3.990 41.840 411.845 47.240 ;
        RECT 4.400 40.440 411.845 41.840 ;
        RECT 3.990 36.400 411.845 40.440 ;
        RECT 3.990 35.000 411.445 36.400 ;
        RECT 3.990 29.600 411.845 35.000 ;
        RECT 4.400 28.200 411.845 29.600 ;
        RECT 3.990 24.160 411.845 28.200 ;
        RECT 3.990 22.760 411.445 24.160 ;
        RECT 3.990 17.360 411.845 22.760 ;
        RECT 4.400 15.960 411.845 17.360 ;
        RECT 3.990 10.715 411.845 15.960 ;
      LAYER met4 ;
        RECT 9.495 12.415 20.640 407.825 ;
        RECT 23.040 12.415 23.940 407.825 ;
        RECT 26.340 12.415 70.640 407.825 ;
        RECT 73.040 12.415 73.940 407.825 ;
        RECT 76.340 12.415 120.640 407.825 ;
        RECT 123.040 12.415 123.940 407.825 ;
        RECT 126.340 12.415 170.640 407.825 ;
        RECT 173.040 12.415 173.940 407.825 ;
        RECT 176.340 12.415 220.640 407.825 ;
        RECT 223.040 12.415 223.940 407.825 ;
        RECT 226.340 12.415 270.640 407.825 ;
        RECT 273.040 12.415 273.940 407.825 ;
        RECT 276.340 12.415 320.640 407.825 ;
        RECT 323.040 12.415 323.940 407.825 ;
        RECT 326.340 12.415 370.640 407.825 ;
        RECT 373.040 12.415 373.940 407.825 ;
        RECT 376.340 12.415 403.585 407.825 ;
  END
END pipelined_mult
END LIBRARY

