module pipelined_mult (clk,
    rst,
    a,
    b,
    p,
    VPWR,
    VGND);
 input clk;
 input rst;
 input [31:0] a;
 input [31:0] b;
 output [63:0] p;
 inout VPWR;
 inout VGND;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire \a_h[0] ;
 wire \a_h[10] ;
 wire \a_h[11] ;
 wire \a_h[12] ;
 wire \a_h[13] ;
 wire \a_h[14] ;
 wire \a_h[15] ;
 wire \a_h[1] ;
 wire \a_h[2] ;
 wire \a_h[3] ;
 wire \a_h[4] ;
 wire \a_h[5] ;
 wire \a_h[6] ;
 wire \a_h[7] ;
 wire \a_h[8] ;
 wire \a_h[9] ;
 wire \a_l[0] ;
 wire \a_l[10] ;
 wire \a_l[11] ;
 wire \a_l[12] ;
 wire \a_l[13] ;
 wire \a_l[14] ;
 wire \a_l[15] ;
 wire \a_l[1] ;
 wire \a_l[2] ;
 wire \a_l[3] ;
 wire \a_l[4] ;
 wire \a_l[5] ;
 wire \a_l[6] ;
 wire \a_l[7] ;
 wire \a_l[8] ;
 wire \a_l[9] ;
 wire \b_h[0] ;
 wire \b_h[10] ;
 wire \b_h[11] ;
 wire \b_h[12] ;
 wire \b_h[13] ;
 wire \b_h[14] ;
 wire \b_h[15] ;
 wire \b_h[1] ;
 wire \b_h[2] ;
 wire \b_h[3] ;
 wire \b_h[4] ;
 wire \b_h[5] ;
 wire \b_h[6] ;
 wire \b_h[7] ;
 wire \b_h[8] ;
 wire \b_h[9] ;
 wire \b_l[0] ;
 wire \b_l[10] ;
 wire \b_l[11] ;
 wire \b_l[12] ;
 wire \b_l[13] ;
 wire \b_l[14] ;
 wire \b_l[15] ;
 wire \b_l[1] ;
 wire \b_l[2] ;
 wire \b_l[3] ;
 wire \b_l[4] ;
 wire \b_l[5] ;
 wire \b_l[6] ;
 wire \b_l[7] ;
 wire \b_l[8] ;
 wire \b_l[9] ;
 wire \mid_sum[0] ;
 wire \mid_sum[10] ;
 wire \mid_sum[11] ;
 wire \mid_sum[12] ;
 wire \mid_sum[13] ;
 wire \mid_sum[14] ;
 wire \mid_sum[15] ;
 wire \mid_sum[16] ;
 wire \mid_sum[17] ;
 wire \mid_sum[18] ;
 wire \mid_sum[19] ;
 wire \mid_sum[1] ;
 wire \mid_sum[20] ;
 wire \mid_sum[21] ;
 wire \mid_sum[22] ;
 wire \mid_sum[23] ;
 wire \mid_sum[24] ;
 wire \mid_sum[25] ;
 wire \mid_sum[26] ;
 wire \mid_sum[27] ;
 wire \mid_sum[28] ;
 wire \mid_sum[29] ;
 wire \mid_sum[2] ;
 wire \mid_sum[30] ;
 wire \mid_sum[31] ;
 wire \mid_sum[32] ;
 wire \mid_sum[3] ;
 wire \mid_sum[4] ;
 wire \mid_sum[5] ;
 wire \mid_sum[6] ;
 wire \mid_sum[7] ;
 wire \mid_sum[8] ;
 wire \mid_sum[9] ;
 wire \p_hh[0] ;
 wire \p_hh[10] ;
 wire \p_hh[11] ;
 wire \p_hh[12] ;
 wire \p_hh[13] ;
 wire \p_hh[14] ;
 wire \p_hh[15] ;
 wire \p_hh[16] ;
 wire \p_hh[17] ;
 wire \p_hh[18] ;
 wire \p_hh[19] ;
 wire \p_hh[1] ;
 wire \p_hh[20] ;
 wire \p_hh[21] ;
 wire \p_hh[22] ;
 wire \p_hh[23] ;
 wire \p_hh[24] ;
 wire \p_hh[25] ;
 wire \p_hh[26] ;
 wire \p_hh[27] ;
 wire \p_hh[28] ;
 wire \p_hh[29] ;
 wire \p_hh[2] ;
 wire \p_hh[30] ;
 wire \p_hh[31] ;
 wire \p_hh[3] ;
 wire \p_hh[4] ;
 wire \p_hh[5] ;
 wire \p_hh[6] ;
 wire \p_hh[7] ;
 wire \p_hh[8] ;
 wire \p_hh[9] ;
 wire \p_hh_pipe[0] ;
 wire \p_hh_pipe[10] ;
 wire \p_hh_pipe[11] ;
 wire \p_hh_pipe[12] ;
 wire \p_hh_pipe[13] ;
 wire \p_hh_pipe[14] ;
 wire \p_hh_pipe[15] ;
 wire \p_hh_pipe[16] ;
 wire \p_hh_pipe[17] ;
 wire \p_hh_pipe[18] ;
 wire \p_hh_pipe[19] ;
 wire \p_hh_pipe[1] ;
 wire \p_hh_pipe[20] ;
 wire \p_hh_pipe[21] ;
 wire \p_hh_pipe[22] ;
 wire \p_hh_pipe[23] ;
 wire \p_hh_pipe[24] ;
 wire \p_hh_pipe[25] ;
 wire \p_hh_pipe[26] ;
 wire \p_hh_pipe[27] ;
 wire \p_hh_pipe[28] ;
 wire \p_hh_pipe[29] ;
 wire \p_hh_pipe[2] ;
 wire \p_hh_pipe[30] ;
 wire \p_hh_pipe[31] ;
 wire \p_hh_pipe[3] ;
 wire \p_hh_pipe[4] ;
 wire \p_hh_pipe[5] ;
 wire \p_hh_pipe[6] ;
 wire \p_hh_pipe[7] ;
 wire \p_hh_pipe[8] ;
 wire \p_hh_pipe[9] ;
 wire \p_hl[0] ;
 wire \p_hl[10] ;
 wire \p_hl[11] ;
 wire \p_hl[12] ;
 wire \p_hl[13] ;
 wire \p_hl[14] ;
 wire \p_hl[15] ;
 wire \p_hl[16] ;
 wire \p_hl[17] ;
 wire \p_hl[18] ;
 wire \p_hl[19] ;
 wire \p_hl[1] ;
 wire \p_hl[20] ;
 wire \p_hl[21] ;
 wire \p_hl[22] ;
 wire \p_hl[23] ;
 wire \p_hl[24] ;
 wire \p_hl[25] ;
 wire \p_hl[26] ;
 wire \p_hl[27] ;
 wire \p_hl[28] ;
 wire \p_hl[29] ;
 wire \p_hl[2] ;
 wire \p_hl[30] ;
 wire \p_hl[31] ;
 wire \p_hl[3] ;
 wire \p_hl[4] ;
 wire \p_hl[5] ;
 wire \p_hl[6] ;
 wire \p_hl[7] ;
 wire \p_hl[8] ;
 wire \p_hl[9] ;
 wire \p_lh[0] ;
 wire \p_lh[10] ;
 wire \p_lh[11] ;
 wire \p_lh[12] ;
 wire \p_lh[13] ;
 wire \p_lh[14] ;
 wire \p_lh[15] ;
 wire \p_lh[16] ;
 wire \p_lh[17] ;
 wire \p_lh[18] ;
 wire \p_lh[19] ;
 wire \p_lh[1] ;
 wire \p_lh[20] ;
 wire \p_lh[21] ;
 wire \p_lh[22] ;
 wire \p_lh[23] ;
 wire \p_lh[24] ;
 wire \p_lh[25] ;
 wire \p_lh[26] ;
 wire \p_lh[27] ;
 wire \p_lh[28] ;
 wire \p_lh[29] ;
 wire \p_lh[2] ;
 wire \p_lh[30] ;
 wire \p_lh[31] ;
 wire \p_lh[3] ;
 wire \p_lh[4] ;
 wire \p_lh[5] ;
 wire \p_lh[6] ;
 wire \p_lh[7] ;
 wire \p_lh[8] ;
 wire \p_lh[9] ;
 wire \p_ll[0] ;
 wire \p_ll[10] ;
 wire \p_ll[11] ;
 wire \p_ll[12] ;
 wire \p_ll[13] ;
 wire \p_ll[14] ;
 wire \p_ll[15] ;
 wire \p_ll[16] ;
 wire \p_ll[17] ;
 wire \p_ll[18] ;
 wire \p_ll[19] ;
 wire \p_ll[1] ;
 wire \p_ll[20] ;
 wire \p_ll[21] ;
 wire \p_ll[22] ;
 wire \p_ll[23] ;
 wire \p_ll[24] ;
 wire \p_ll[25] ;
 wire \p_ll[26] ;
 wire \p_ll[27] ;
 wire \p_ll[28] ;
 wire \p_ll[29] ;
 wire \p_ll[2] ;
 wire \p_ll[30] ;
 wire \p_ll[31] ;
 wire \p_ll[3] ;
 wire \p_ll[4] ;
 wire \p_ll[5] ;
 wire \p_ll[6] ;
 wire \p_ll[7] ;
 wire \p_ll[8] ;
 wire \p_ll[9] ;
 wire \p_ll_pipe[0] ;
 wire \p_ll_pipe[10] ;
 wire \p_ll_pipe[11] ;
 wire \p_ll_pipe[12] ;
 wire \p_ll_pipe[13] ;
 wire \p_ll_pipe[14] ;
 wire \p_ll_pipe[15] ;
 wire \p_ll_pipe[16] ;
 wire \p_ll_pipe[17] ;
 wire \p_ll_pipe[18] ;
 wire \p_ll_pipe[19] ;
 wire \p_ll_pipe[1] ;
 wire \p_ll_pipe[20] ;
 wire \p_ll_pipe[21] ;
 wire \p_ll_pipe[22] ;
 wire \p_ll_pipe[23] ;
 wire \p_ll_pipe[24] ;
 wire \p_ll_pipe[25] ;
 wire \p_ll_pipe[26] ;
 wire \p_ll_pipe[27] ;
 wire \p_ll_pipe[28] ;
 wire \p_ll_pipe[29] ;
 wire \p_ll_pipe[2] ;
 wire \p_ll_pipe[30] ;
 wire \p_ll_pipe[31] ;
 wire \p_ll_pipe[3] ;
 wire \p_ll_pipe[4] ;
 wire \p_ll_pipe[5] ;
 wire \p_ll_pipe[6] ;
 wire \p_ll_pipe[7] ;
 wire \p_ll_pipe[8] ;
 wire \p_ll_pipe[9] ;
 wire \term_high[32] ;
 wire \term_high[33] ;
 wire \term_high[34] ;
 wire \term_high[35] ;
 wire \term_high[36] ;
 wire \term_high[37] ;
 wire \term_high[38] ;
 wire \term_high[39] ;
 wire \term_high[40] ;
 wire \term_high[41] ;
 wire \term_high[42] ;
 wire \term_high[43] ;
 wire \term_high[44] ;
 wire \term_high[45] ;
 wire \term_high[46] ;
 wire \term_high[47] ;
 wire \term_high[48] ;
 wire \term_high[49] ;
 wire \term_high[50] ;
 wire \term_high[51] ;
 wire \term_high[52] ;
 wire \term_high[53] ;
 wire \term_high[54] ;
 wire \term_high[55] ;
 wire \term_high[56] ;
 wire \term_high[57] ;
 wire \term_high[58] ;
 wire \term_high[59] ;
 wire \term_high[60] ;
 wire \term_high[61] ;
 wire \term_high[62] ;
 wire \term_high[63] ;
 wire \term_low[0] ;
 wire \term_low[10] ;
 wire \term_low[11] ;
 wire \term_low[12] ;
 wire \term_low[13] ;
 wire \term_low[14] ;
 wire \term_low[15] ;
 wire \term_low[16] ;
 wire \term_low[17] ;
 wire \term_low[18] ;
 wire \term_low[19] ;
 wire \term_low[1] ;
 wire \term_low[20] ;
 wire \term_low[21] ;
 wire \term_low[22] ;
 wire \term_low[23] ;
 wire \term_low[24] ;
 wire \term_low[25] ;
 wire \term_low[26] ;
 wire \term_low[27] ;
 wire \term_low[28] ;
 wire \term_low[29] ;
 wire \term_low[2] ;
 wire \term_low[30] ;
 wire \term_low[31] ;
 wire \term_low[3] ;
 wire \term_low[4] ;
 wire \term_low[5] ;
 wire \term_low[6] ;
 wire \term_low[7] ;
 wire \term_low[8] ;
 wire \term_low[9] ;
 wire \term_mid[16] ;
 wire \term_mid[17] ;
 wire \term_mid[18] ;
 wire \term_mid[19] ;
 wire \term_mid[20] ;
 wire \term_mid[21] ;
 wire \term_mid[22] ;
 wire \term_mid[23] ;
 wire \term_mid[24] ;
 wire \term_mid[25] ;
 wire \term_mid[26] ;
 wire \term_mid[27] ;
 wire \term_mid[28] ;
 wire \term_mid[29] ;
 wire \term_mid[30] ;
 wire \term_mid[31] ;
 wire \term_mid[32] ;
 wire \term_mid[33] ;
 wire \term_mid[34] ;
 wire \term_mid[35] ;
 wire \term_mid[36] ;
 wire \term_mid[37] ;
 wire \term_mid[38] ;
 wire \term_mid[39] ;
 wire \term_mid[40] ;
 wire \term_mid[41] ;
 wire \term_mid[42] ;
 wire \term_mid[43] ;
 wire \term_mid[44] ;
 wire \term_mid[45] ;
 wire \term_mid[46] ;
 wire \term_mid[47] ;
 wire \term_mid[48] ;

 sky130_fd_sc_hd__inv_2 _10180_ (.A(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09144_));
 sky130_fd_sc_hd__inv_2 _10181_ (.A(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_2 _10182_ (.A(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09166_));
 sky130_fd_sc_hd__inv_2 _10183_ (.A(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09177_));
 sky130_fd_sc_hd__inv_2 _10184_ (.A(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09188_));
 sky130_fd_sc_hd__inv_2 _10185_ (.A(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09199_));
 sky130_fd_sc_hd__inv_2 _10186_ (.A(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09210_));
 sky130_fd_sc_hd__inv_2 _10187_ (.A(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09220_));
 sky130_fd_sc_hd__inv_2 _10188_ (.A(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09231_));
 sky130_fd_sc_hd__inv_2 _10189_ (.A(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09242_));
 sky130_fd_sc_hd__inv_2 _10190_ (.A(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09253_));
 sky130_fd_sc_hd__inv_2 _10191_ (.A(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09264_));
 sky130_fd_sc_hd__inv_2 _10192_ (.A(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09275_));
 sky130_fd_sc_hd__inv_2 _10193_ (.A(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09286_));
 sky130_fd_sc_hd__inv_2 _10194_ (.A(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09297_));
 sky130_fd_sc_hd__inv_2 _10195_ (.A(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09308_));
 sky130_fd_sc_hd__inv_2 _10196_ (.A(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09319_));
 sky130_fd_sc_hd__inv_2 _10197_ (.A(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09329_));
 sky130_fd_sc_hd__inv_2 _10198_ (.A(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09340_));
 sky130_fd_sc_hd__inv_2 _10199_ (.A(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09351_));
 sky130_fd_sc_hd__inv_2 _10200_ (.A(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09362_));
 sky130_fd_sc_hd__inv_2 _10201_ (.A(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09373_));
 sky130_fd_sc_hd__inv_2 _10202_ (.A(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09384_));
 sky130_fd_sc_hd__inv_2 _10203_ (.A(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09395_));
 sky130_fd_sc_hd__inv_2 _10204_ (.A(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09406_));
 sky130_fd_sc_hd__inv_2 _10205_ (.A(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09417_));
 sky130_fd_sc_hd__inv_2 _10206_ (.A(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09428_));
 sky130_fd_sc_hd__inv_2 _10207_ (.A(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09439_));
 sky130_fd_sc_hd__inv_2 _10208_ (.A(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09449_));
 sky130_fd_sc_hd__inv_2 _10209_ (.A(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09460_));
 sky130_fd_sc_hd__inv_2 _10210_ (.A(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09471_));
 sky130_fd_sc_hd__inv_2 _10211_ (.A(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09482_));
 sky130_fd_sc_hd__inv_2 _10212_ (.A(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09493_));
 sky130_fd_sc_hd__inv_2 _10213_ (.A(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09504_));
 sky130_fd_sc_hd__inv_2 _10214_ (.A(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09515_));
 sky130_fd_sc_hd__inv_2 _10215_ (.A(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09526_));
 sky130_fd_sc_hd__inv_2 _10216_ (.A(\p_hl[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09537_));
 sky130_fd_sc_hd__inv_2 _10217_ (.A(\p_lh[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09548_));
 sky130_fd_sc_hd__inv_2 _10218_ (.A(\p_hl[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09559_));
 sky130_fd_sc_hd__inv_2 _10219_ (.A(\p_lh[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09570_));
 sky130_fd_sc_hd__inv_2 _10220_ (.A(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09581_));
 sky130_fd_sc_hd__inv_2 _10221_ (.A(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09592_));
 sky130_fd_sc_hd__inv_2 _10222_ (.A(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09602_));
 sky130_fd_sc_hd__inv_2 _10223_ (.A(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09613_));
 sky130_fd_sc_hd__inv_2 _10224_ (.A(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09624_));
 sky130_fd_sc_hd__inv_2 _10225_ (.A(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09635_));
 sky130_fd_sc_hd__inv_2 _10226_ (.A(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09646_));
 sky130_fd_sc_hd__inv_2 _10227_ (.A(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09657_));
 sky130_fd_sc_hd__inv_2 _10228_ (.A(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09668_));
 sky130_fd_sc_hd__inv_2 _10229_ (.A(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09679_));
 sky130_fd_sc_hd__inv_2 _10230_ (.A(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09690_));
 sky130_fd_sc_hd__and2_2 _10231_ (.A(_09690_),
    .B(b[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00000_));
 sky130_fd_sc_hd__and2_2 _10232_ (.A(_09690_),
    .B(b[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00001_));
 sky130_fd_sc_hd__and2_2 _10233_ (.A(_09690_),
    .B(b[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00002_));
 sky130_fd_sc_hd__and2_2 _10234_ (.A(_09690_),
    .B(b[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00003_));
 sky130_fd_sc_hd__and2_2 _10235_ (.A(_09690_),
    .B(b[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00004_));
 sky130_fd_sc_hd__and2_2 _10236_ (.A(_09690_),
    .B(b[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00005_));
 sky130_fd_sc_hd__and2_2 _10237_ (.A(_09690_),
    .B(b[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00006_));
 sky130_fd_sc_hd__and2_2 _10238_ (.A(_09690_),
    .B(b[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00007_));
 sky130_fd_sc_hd__and2_2 _10239_ (.A(_09690_),
    .B(b[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00008_));
 sky130_fd_sc_hd__and2_2 _10240_ (.A(_09690_),
    .B(b[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00009_));
 sky130_fd_sc_hd__and2_2 _10241_ (.A(_09690_),
    .B(b[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00010_));
 sky130_fd_sc_hd__and2_2 _10242_ (.A(_09690_),
    .B(b[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00011_));
 sky130_fd_sc_hd__and2_2 _10243_ (.A(_09690_),
    .B(b[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00012_));
 sky130_fd_sc_hd__and2_2 _10244_ (.A(_09690_),
    .B(b[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00013_));
 sky130_fd_sc_hd__and2_2 _10245_ (.A(_09690_),
    .B(b[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00014_));
 sky130_fd_sc_hd__and2_2 _10246_ (.A(_09690_),
    .B(b[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00015_));
 sky130_fd_sc_hd__and2_2 _10247_ (.A(_09690_),
    .B(\term_low[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00016_));
 sky130_fd_sc_hd__and2_2 _10248_ (.A(_09690_),
    .B(\term_low[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00017_));
 sky130_fd_sc_hd__and2_2 _10249_ (.A(_09690_),
    .B(\term_low[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00018_));
 sky130_fd_sc_hd__and2_2 _10250_ (.A(_09690_),
    .B(\term_low[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00019_));
 sky130_fd_sc_hd__and2_2 _10251_ (.A(_09690_),
    .B(\term_low[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00020_));
 sky130_fd_sc_hd__and2_2 _10252_ (.A(_09690_),
    .B(\term_low[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00021_));
 sky130_fd_sc_hd__and2_2 _10253_ (.A(_09690_),
    .B(\term_low[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00022_));
 sky130_fd_sc_hd__and2_2 _10254_ (.A(_09690_),
    .B(\term_low[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00023_));
 sky130_fd_sc_hd__and2_2 _10255_ (.A(_09690_),
    .B(\term_low[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00024_));
 sky130_fd_sc_hd__and2_2 _10256_ (.A(_09690_),
    .B(\term_low[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00025_));
 sky130_fd_sc_hd__and2_2 _10257_ (.A(_09690_),
    .B(\term_low[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00026_));
 sky130_fd_sc_hd__and2_2 _10258_ (.A(_09690_),
    .B(\term_low[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00027_));
 sky130_fd_sc_hd__and2_2 _10259_ (.A(_09690_),
    .B(\term_low[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00028_));
 sky130_fd_sc_hd__and2_2 _10260_ (.A(_09690_),
    .B(\term_low[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00029_));
 sky130_fd_sc_hd__and2_2 _10261_ (.A(_09690_),
    .B(\term_low[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00030_));
 sky130_fd_sc_hd__and2_2 _10262_ (.A(_09690_),
    .B(\term_low[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_2 _10263_ (.A(\term_low[16] ),
    .B(\term_mid[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10018_));
 sky130_fd_sc_hd__a21oi_2 _10264_ (.A1(\term_low[16] ),
    .A2(\term_mid[16] ),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10029_));
 sky130_fd_sc_hd__o21a_2 _10265_ (.A1(\term_low[16] ),
    .A2(\term_mid[16] ),
    .B1(_10029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00032_));
 sky130_fd_sc_hd__and2_2 _10266_ (.A(\term_low[17] ),
    .B(\term_mid[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10050_));
 sky130_fd_sc_hd__nand2_2 _10267_ (.A(\term_low[17] ),
    .B(\term_mid[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10061_));
 sky130_fd_sc_hd__nor2_2 _10268_ (.A(\term_low[17] ),
    .B(\term_mid[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10072_));
 sky130_fd_sc_hd__or2_2 _10269_ (.A(_10018_),
    .B(_10072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10083_));
 sky130_fd_sc_hd__a2bb2o_2 _10270_ (.A1_N(_10050_),
    .A2_N(_10072_),
    .B1(\term_low[16] ),
    .B2(\term_mid[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10094_));
 sky130_fd_sc_hd__o211a_2 _10271_ (.A1(_10083_),
    .A2(_10050_),
    .B1(_09690_),
    .C1(_10094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00033_));
 sky130_fd_sc_hd__o21ai_2 _10272_ (.A1(_10018_),
    .A2(_10072_),
    .B1(_10061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10115_));
 sky130_fd_sc_hd__nor2_2 _10273_ (.A(\term_low[18] ),
    .B(\term_mid[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10126_));
 sky130_fd_sc_hd__and2_2 _10274_ (.A(\term_low[18] ),
    .B(\term_mid[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10137_));
 sky130_fd_sc_hd__nand2_2 _10275_ (.A(\term_low[18] ),
    .B(\term_mid[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10148_));
 sky130_fd_sc_hd__nor2_2 _10276_ (.A(_10126_),
    .B(_10137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10158_));
 sky130_fd_sc_hd__nand2_2 _10277_ (.A(_10158_),
    .B(_10115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10169_));
 sky130_fd_sc_hd__a21oi_2 _10278_ (.A1(_10158_),
    .A2(_10115_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00450_));
 sky130_fd_sc_hd__o21a_2 _10279_ (.A1(_10115_),
    .A2(_10158_),
    .B1(_00450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00034_));
 sky130_fd_sc_hd__or2_2 _10280_ (.A(\term_low[19] ),
    .B(\term_mid[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00471_));
 sky130_fd_sc_hd__nand2_2 _10281_ (.A(\term_low[19] ),
    .B(\term_mid[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_2 _10282_ (.A(_00471_),
    .B(_00482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00493_));
 sky130_fd_sc_hd__a21oi_2 _10283_ (.A1(_10148_),
    .A2(_10169_),
    .B1(_00493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00504_));
 sky130_fd_sc_hd__a31o_2 _10284_ (.A1(_10148_),
    .A2(_10169_),
    .A3(_00493_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_2 _10285_ (.A(_00504_),
    .B(_00515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00035_));
 sky130_fd_sc_hd__nand2_2 _10286_ (.A(\term_low[20] ),
    .B(\term_mid[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00536_));
 sky130_fd_sc_hd__nand3_2 _10287_ (.A(_10148_),
    .B(_10169_),
    .C(_00482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00547_));
 sky130_fd_sc_hd__o21ai_2 _10288_ (.A1(\term_low[19] ),
    .A2(\term_mid[19] ),
    .B1(_00547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00558_));
 sky130_fd_sc_hd__o211ai_2 _10289_ (.A1(\term_low[20] ),
    .A2(\term_mid[20] ),
    .B1(_00471_),
    .C1(_00547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00569_));
 sky130_fd_sc_hd__xnor2_2 _10290_ (.A(\term_low[20] ),
    .B(\term_mid[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00579_));
 sky130_fd_sc_hd__a21oi_2 _10291_ (.A1(_00558_),
    .A2(_00579_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00590_));
 sky130_fd_sc_hd__o21a_2 _10292_ (.A1(_00558_),
    .A2(_00579_),
    .B1(_00590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00036_));
 sky130_fd_sc_hd__nor2_2 _10293_ (.A(\term_low[21] ),
    .B(\term_mid[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00611_));
 sky130_fd_sc_hd__and2_2 _10294_ (.A(\term_low[21] ),
    .B(\term_mid[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00622_));
 sky130_fd_sc_hd__nand2_2 _10295_ (.A(\term_low[21] ),
    .B(\term_mid[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00633_));
 sky130_fd_sc_hd__a211o_2 _10296_ (.A1(_00536_),
    .A2(_00569_),
    .B1(_00611_),
    .C1(_00622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00644_));
 sky130_fd_sc_hd__o211ai_2 _10297_ (.A1(_00611_),
    .A2(_00622_),
    .B1(_00536_),
    .C1(_00569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00655_));
 sky130_fd_sc_hd__and3_2 _10298_ (.A(_09690_),
    .B(_00644_),
    .C(_00655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00037_));
 sky130_fd_sc_hd__nor2_2 _10299_ (.A(\term_low[22] ),
    .B(\term_mid[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00676_));
 sky130_fd_sc_hd__or2_2 _10300_ (.A(\term_low[22] ),
    .B(\term_mid[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00687_));
 sky130_fd_sc_hd__nand2_2 _10301_ (.A(\term_low[22] ),
    .B(\term_mid[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_2 _10302_ (.A(_00687_),
    .B(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00709_));
 sky130_fd_sc_hd__nand3_2 _10303_ (.A(_00536_),
    .B(_00569_),
    .C(_00633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00719_));
 sky130_fd_sc_hd__o21ai_2 _10304_ (.A1(\term_low[21] ),
    .A2(\term_mid[21] ),
    .B1(_00719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00730_));
 sky130_fd_sc_hd__a21oi_2 _10305_ (.A1(_00709_),
    .A2(_00730_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00741_));
 sky130_fd_sc_hd__o21a_2 _10306_ (.A1(_00709_),
    .A2(_00730_),
    .B1(_00741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00038_));
 sky130_fd_sc_hd__o211ai_2 _10307_ (.A1(\term_low[21] ),
    .A2(\term_mid[21] ),
    .B1(_00687_),
    .C1(_00719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00762_));
 sky130_fd_sc_hd__o21ai_2 _10308_ (.A1(_00676_),
    .A2(_00730_),
    .B1(_00698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00773_));
 sky130_fd_sc_hd__nand2_2 _10309_ (.A(\term_low[23] ),
    .B(\term_mid[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00784_));
 sky130_fd_sc_hd__or2_2 _10310_ (.A(\term_low[23] ),
    .B(\term_mid[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00795_));
 sky130_fd_sc_hd__a21oi_2 _10311_ (.A1(_00784_),
    .A2(_00795_),
    .B1(_00773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00806_));
 sky130_fd_sc_hd__a311oi_2 _10312_ (.A1(_00773_),
    .A2(_00784_),
    .A3(_00795_),
    .B1(_00806_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00039_));
 sky130_fd_sc_hd__xor2_2 _10313_ (.A(\term_low[24] ),
    .B(\term_mid[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00827_));
 sky130_fd_sc_hd__nand3_2 _10314_ (.A(_00698_),
    .B(_00762_),
    .C(_00784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00838_));
 sky130_fd_sc_hd__a21o_2 _10315_ (.A1(_00795_),
    .A2(_00838_),
    .B1(_00827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00849_));
 sky130_fd_sc_hd__and3_2 _10316_ (.A(_00795_),
    .B(_00838_),
    .C(_00827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00859_));
 sky130_fd_sc_hd__o211ai_2 _10317_ (.A1(\term_low[23] ),
    .A2(\term_mid[23] ),
    .B1(_00827_),
    .C1(_00838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00870_));
 sky130_fd_sc_hd__and3_2 _10318_ (.A(_09690_),
    .B(_00849_),
    .C(_00870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00040_));
 sky130_fd_sc_hd__nor2_2 _10319_ (.A(\term_low[25] ),
    .B(\term_mid[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00891_));
 sky130_fd_sc_hd__and2_2 _10320_ (.A(\term_low[25] ),
    .B(\term_mid[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00902_));
 sky130_fd_sc_hd__nor2_2 _10321_ (.A(_00891_),
    .B(_00902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00913_));
 sky130_fd_sc_hd__a21o_2 _10322_ (.A1(\term_low[24] ),
    .A2(\term_mid[24] ),
    .B1(_00859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00924_));
 sky130_fd_sc_hd__o21ai_2 _10323_ (.A1(_00913_),
    .A2(_00924_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00935_));
 sky130_fd_sc_hd__a21oi_2 _10324_ (.A1(_00913_),
    .A2(_00924_),
    .B1(_00935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00041_));
 sky130_fd_sc_hd__and2_2 _10325_ (.A(\term_low[26] ),
    .B(\term_mid[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00956_));
 sky130_fd_sc_hd__nor2_2 _10326_ (.A(\term_low[26] ),
    .B(\term_mid[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00967_));
 sky130_fd_sc_hd__a21oi_2 _10327_ (.A1(\term_low[24] ),
    .A2(\term_mid[24] ),
    .B1(_00902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_2 _10328_ (.A(_00870_),
    .B(_00978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00988_));
 sky130_fd_sc_hd__a2bb2o_2 _10329_ (.A1_N(\term_low[25] ),
    .A2_N(\term_mid[25] ),
    .B1(_00978_),
    .B2(_00870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00999_));
 sky130_fd_sc_hd__o21ai_2 _10330_ (.A1(_00956_),
    .A2(_00967_),
    .B1(_00999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01010_));
 sky130_fd_sc_hd__or3_2 _10331_ (.A(_00956_),
    .B(_00967_),
    .C(_00999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01021_));
 sky130_fd_sc_hd__and3_2 _10332_ (.A(_09690_),
    .B(_01010_),
    .C(_01021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00042_));
 sky130_fd_sc_hd__xor2_2 _10333_ (.A(\term_low[27] ),
    .B(\term_mid[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01042_));
 sky130_fd_sc_hd__a21bo_2 _10334_ (.A1(\term_low[26] ),
    .A2(\term_mid[26] ),
    .B1_N(_01021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01053_));
 sky130_fd_sc_hd__a21oi_2 _10335_ (.A1(_01053_),
    .A2(_01042_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01064_));
 sky130_fd_sc_hd__o21a_2 _10336_ (.A1(_01042_),
    .A2(_01053_),
    .B1(_01064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00043_));
 sky130_fd_sc_hd__nor2_2 _10337_ (.A(\term_low[28] ),
    .B(\term_mid[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01084_));
 sky130_fd_sc_hd__and2_2 _10338_ (.A(\term_low[28] ),
    .B(\term_mid[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01095_));
 sky130_fd_sc_hd__or2_2 _10339_ (.A(_01084_),
    .B(_01095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01106_));
 sky130_fd_sc_hd__o211a_2 _10340_ (.A1(\term_low[27] ),
    .A2(\term_mid[27] ),
    .B1(\term_low[26] ),
    .C1(\term_mid[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01117_));
 sky130_fd_sc_hd__a21o_2 _10341_ (.A1(\term_low[27] ),
    .A2(\term_mid[27] ),
    .B1(_01117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01128_));
 sky130_fd_sc_hd__or4b_2 _10342_ (.A(_00891_),
    .B(_00956_),
    .C(_00967_),
    .D_N(_01042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01139_));
 sky130_fd_sc_hd__inv_2 _10343_ (.A(_01139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01150_));
 sky130_fd_sc_hd__a21oi_2 _10344_ (.A1(_00988_),
    .A2(_01150_),
    .B1(_01128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01161_));
 sky130_fd_sc_hd__o21ai_2 _10345_ (.A1(_01106_),
    .A2(_01161_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01172_));
 sky130_fd_sc_hd__a21oi_2 _10346_ (.A1(_01106_),
    .A2(_01161_),
    .B1(_01172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00044_));
 sky130_fd_sc_hd__and2_2 _10347_ (.A(\term_low[29] ),
    .B(\term_mid[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01192_));
 sky130_fd_sc_hd__nor2_2 _10348_ (.A(\term_low[29] ),
    .B(\term_mid[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01203_));
 sky130_fd_sc_hd__nor2_2 _10349_ (.A(_01192_),
    .B(_01203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01214_));
 sky130_fd_sc_hd__o21bai_2 _10350_ (.A1(_01106_),
    .A2(_01161_),
    .B1_N(_01095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01225_));
 sky130_fd_sc_hd__a21oi_2 _10351_ (.A1(_01225_),
    .A2(_01214_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01236_));
 sky130_fd_sc_hd__o21a_2 _10352_ (.A1(_01214_),
    .A2(_01225_),
    .B1(_01236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00045_));
 sky130_fd_sc_hd__nand2_2 _10353_ (.A(\term_low[30] ),
    .B(\term_mid[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01257_));
 sky130_fd_sc_hd__xnor2_2 _10354_ (.A(\term_low[30] ),
    .B(\term_mid[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01268_));
 sky130_fd_sc_hd__o211a_2 _10355_ (.A1(\term_low[29] ),
    .A2(\term_mid[29] ),
    .B1(\term_low[28] ),
    .C1(\term_mid[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01278_));
 sky130_fd_sc_hd__a21oi_2 _10356_ (.A1(\term_low[29] ),
    .A2(\term_mid[29] ),
    .B1(_01278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01289_));
 sky130_fd_sc_hd__or4_2 _10357_ (.A(_01084_),
    .B(_01095_),
    .C(_01192_),
    .D(_01203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01300_));
 sky130_fd_sc_hd__o21ai_2 _10358_ (.A1(_01161_),
    .A2(_01300_),
    .B1(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01311_));
 sky130_fd_sc_hd__o21a_2 _10359_ (.A1(_01161_),
    .A2(_01300_),
    .B1(_01289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01322_));
 sky130_fd_sc_hd__o21ai_2 _10360_ (.A1(_01268_),
    .A2(_01322_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01333_));
 sky130_fd_sc_hd__a21oi_2 _10361_ (.A1(_01268_),
    .A2(_01322_),
    .B1(_01333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00046_));
 sky130_fd_sc_hd__nor2_2 _10362_ (.A(\term_low[31] ),
    .B(\term_mid[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01354_));
 sky130_fd_sc_hd__and2_2 _10363_ (.A(\term_low[31] ),
    .B(\term_mid[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01364_));
 sky130_fd_sc_hd__nor2_2 _10364_ (.A(_01354_),
    .B(_01364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01375_));
 sky130_fd_sc_hd__o21ai_2 _10365_ (.A1(_01268_),
    .A2(_01322_),
    .B1(_01257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01386_));
 sky130_fd_sc_hd__a21oi_2 _10366_ (.A1(_01386_),
    .A2(_01375_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01397_));
 sky130_fd_sc_hd__o21a_2 _10367_ (.A1(_01375_),
    .A2(_01386_),
    .B1(_01397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00047_));
 sky130_fd_sc_hd__xor2_2 _10368_ (.A(\term_mid[32] ),
    .B(\term_high[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01417_));
 sky130_fd_sc_hd__o211a_2 _10369_ (.A1(\term_low[31] ),
    .A2(\term_mid[31] ),
    .B1(\term_low[30] ),
    .C1(\term_mid[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01428_));
 sky130_fd_sc_hd__a21o_2 _10370_ (.A1(\term_low[31] ),
    .A2(\term_mid[31] ),
    .B1(_01428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01439_));
 sky130_fd_sc_hd__nor3_2 _10371_ (.A(_01354_),
    .B(_01364_),
    .C(_01268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01450_));
 sky130_fd_sc_hd__a211o_2 _10372_ (.A1(_01311_),
    .A2(_01450_),
    .B1(_01428_),
    .C1(_01364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01460_));
 sky130_fd_sc_hd__a21oi_2 _10373_ (.A1(_01311_),
    .A2(_01450_),
    .B1(_01439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01471_));
 sky130_fd_sc_hd__and2_2 _10374_ (.A(_01417_),
    .B(_01460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01482_));
 sky130_fd_sc_hd__a21oi_2 _10375_ (.A1(_01417_),
    .A2(_01460_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01493_));
 sky130_fd_sc_hd__o21a_2 _10376_ (.A1(_01417_),
    .A2(_01460_),
    .B1(_01493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00048_));
 sky130_fd_sc_hd__xor2_2 _10377_ (.A(\term_mid[33] ),
    .B(\term_high[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01513_));
 sky130_fd_sc_hd__a21o_2 _10378_ (.A1(\term_mid[32] ),
    .A2(\term_high[32] ),
    .B1(_01482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01524_));
 sky130_fd_sc_hd__a21oi_2 _10379_ (.A1(_01524_),
    .A2(_01513_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01534_));
 sky130_fd_sc_hd__o21a_2 _10380_ (.A1(_01513_),
    .A2(_01524_),
    .B1(_01534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00049_));
 sky130_fd_sc_hd__xor2_2 _10381_ (.A(\term_mid[34] ),
    .B(\term_high[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01554_));
 sky130_fd_sc_hd__a22o_2 _10382_ (.A1(\term_mid[32] ),
    .A2(\term_high[32] ),
    .B1(\term_mid[33] ),
    .B2(\term_high[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01557_));
 sky130_fd_sc_hd__o21a_2 _10383_ (.A1(\term_mid[33] ),
    .A2(\term_high[33] ),
    .B1(_01557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01558_));
 sky130_fd_sc_hd__a31o_2 _10384_ (.A1(_01417_),
    .A2(_01460_),
    .A3(_01513_),
    .B1(_01558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01559_));
 sky130_fd_sc_hd__o221a_2 _10385_ (.A1(\term_mid[33] ),
    .A2(\term_high[33] ),
    .B1(_01557_),
    .B2(_01482_),
    .C1(_01554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01560_));
 sky130_fd_sc_hd__a21oi_2 _10386_ (.A1(_01554_),
    .A2(_01559_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01561_));
 sky130_fd_sc_hd__o21a_2 _10387_ (.A1(_01554_),
    .A2(_01559_),
    .B1(_01561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00050_));
 sky130_fd_sc_hd__xor2_2 _10388_ (.A(\term_mid[35] ),
    .B(\term_high[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01562_));
 sky130_fd_sc_hd__a21o_2 _10389_ (.A1(\term_mid[34] ),
    .A2(\term_high[34] ),
    .B1(_01560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01563_));
 sky130_fd_sc_hd__a21oi_2 _10390_ (.A1(_01563_),
    .A2(_01562_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01564_));
 sky130_fd_sc_hd__o21a_2 _10391_ (.A1(_01562_),
    .A2(_01563_),
    .B1(_01564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00051_));
 sky130_fd_sc_hd__xor2_2 _10392_ (.A(\term_mid[36] ),
    .B(\term_high[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01565_));
 sky130_fd_sc_hd__nand4_2 _10393_ (.A(_01417_),
    .B(_01513_),
    .C(_01554_),
    .D(_01562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01566_));
 sky130_fd_sc_hd__o211a_2 _10394_ (.A1(\term_mid[35] ),
    .A2(\term_high[35] ),
    .B1(\term_mid[34] ),
    .C1(\term_high[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01567_));
 sky130_fd_sc_hd__a21o_2 _10395_ (.A1(\term_mid[35] ),
    .A2(\term_high[35] ),
    .B1(_01567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01568_));
 sky130_fd_sc_hd__a31oi_2 _10396_ (.A1(_01554_),
    .A2(_01558_),
    .A3(_01562_),
    .B1(_01568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01569_));
 sky130_fd_sc_hd__o21ai_2 _10397_ (.A1(_01471_),
    .A2(_01566_),
    .B1(_01569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01570_));
 sky130_fd_sc_hd__or2_2 _10398_ (.A(_01565_),
    .B(_01570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01571_));
 sky130_fd_sc_hd__nand2_2 _10399_ (.A(_01570_),
    .B(_01565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01572_));
 sky130_fd_sc_hd__and3_2 _10400_ (.A(_09690_),
    .B(_01571_),
    .C(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00052_));
 sky130_fd_sc_hd__nor2_2 _10401_ (.A(\term_mid[37] ),
    .B(\term_high[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01573_));
 sky130_fd_sc_hd__and2_2 _10402_ (.A(\term_mid[37] ),
    .B(\term_high[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01574_));
 sky130_fd_sc_hd__nor2_2 _10403_ (.A(_01573_),
    .B(_01574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01575_));
 sky130_fd_sc_hd__a21bo_2 _10404_ (.A1(\term_mid[36] ),
    .A2(\term_high[36] ),
    .B1_N(_01572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01576_));
 sky130_fd_sc_hd__o21a_2 _10405_ (.A1(_01575_),
    .A2(_01576_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01577_));
 sky130_fd_sc_hd__a21boi_2 _10406_ (.A1(_01575_),
    .A2(_01576_),
    .B1_N(_01577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00053_));
 sky130_fd_sc_hd__nor2_2 _10407_ (.A(\term_mid[38] ),
    .B(\term_high[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01578_));
 sky130_fd_sc_hd__and2_2 _10408_ (.A(\term_mid[38] ),
    .B(\term_high[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01579_));
 sky130_fd_sc_hd__nor2_2 _10409_ (.A(_01578_),
    .B(_01579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01580_));
 sky130_fd_sc_hd__and3_2 _10410_ (.A(_01570_),
    .B(_01575_),
    .C(_01565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01581_));
 sky130_fd_sc_hd__o211a_2 _10411_ (.A1(\term_mid[37] ),
    .A2(\term_high[37] ),
    .B1(\term_mid[36] ),
    .C1(\term_high[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01582_));
 sky130_fd_sc_hd__o31a_2 _10412_ (.A1(_01574_),
    .A2(_01581_),
    .A3(_01582_),
    .B1(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01583_));
 sky130_fd_sc_hd__nor2_2 _10413_ (.A(rst),
    .B(_01583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01584_));
 sky130_fd_sc_hd__o41a_2 _10414_ (.A1(_01574_),
    .A2(_01580_),
    .A3(_01581_),
    .A4(_01582_),
    .B1(_01584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00054_));
 sky130_fd_sc_hd__xor2_2 _10415_ (.A(\term_mid[39] ),
    .B(\term_high[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01585_));
 sky130_fd_sc_hd__o21ai_2 _10416_ (.A1(_01579_),
    .A2(_01583_),
    .B1(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01586_));
 sky130_fd_sc_hd__or3_2 _10417_ (.A(_01579_),
    .B(_01583_),
    .C(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01587_));
 sky130_fd_sc_hd__and3_2 _10418_ (.A(_09690_),
    .B(_01586_),
    .C(_01587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00055_));
 sky130_fd_sc_hd__nor2_2 _10419_ (.A(\term_mid[40] ),
    .B(\term_high[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01588_));
 sky130_fd_sc_hd__and2_2 _10420_ (.A(\term_mid[40] ),
    .B(\term_high[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01589_));
 sky130_fd_sc_hd__nor2_2 _10421_ (.A(_01588_),
    .B(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01590_));
 sky130_fd_sc_hd__and4_2 _10422_ (.A(_01565_),
    .B(_01575_),
    .C(_01580_),
    .D(_01585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01591_));
 sky130_fd_sc_hd__o211a_2 _10423_ (.A1(_01574_),
    .A2(_01582_),
    .B1(_01585_),
    .C1(_01580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01592_));
 sky130_fd_sc_hd__o211a_2 _10424_ (.A1(\term_mid[39] ),
    .A2(\term_high[39] ),
    .B1(\term_mid[38] ),
    .C1(\term_high[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01593_));
 sky130_fd_sc_hd__a211o_2 _10425_ (.A1(\term_mid[39] ),
    .A2(\term_high[39] ),
    .B1(_01592_),
    .C1(_01593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01594_));
 sky130_fd_sc_hd__a21o_2 _10426_ (.A1(_01570_),
    .A2(_01591_),
    .B1(_01594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01595_));
 sky130_fd_sc_hd__a21oi_2 _10427_ (.A1(_01595_),
    .A2(_01590_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01596_));
 sky130_fd_sc_hd__o21a_2 _10428_ (.A1(_01590_),
    .A2(_01595_),
    .B1(_01596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00056_));
 sky130_fd_sc_hd__nor2_2 _10429_ (.A(\term_mid[41] ),
    .B(\term_high[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01597_));
 sky130_fd_sc_hd__and2_2 _10430_ (.A(\term_mid[41] ),
    .B(\term_high[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01598_));
 sky130_fd_sc_hd__nor2_2 _10431_ (.A(_01597_),
    .B(_01598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01599_));
 sky130_fd_sc_hd__a21oi_2 _10432_ (.A1(_01595_),
    .A2(_01590_),
    .B1(_01589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01600_));
 sky130_fd_sc_hd__o21a_2 _10433_ (.A1(_01597_),
    .A2(_01598_),
    .B1(_01600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01601_));
 sky130_fd_sc_hd__nor2_2 _10434_ (.A(rst),
    .B(_01601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01602_));
 sky130_fd_sc_hd__o31a_2 _10435_ (.A1(_01597_),
    .A2(_01598_),
    .A3(_01600_),
    .B1(_01602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00057_));
 sky130_fd_sc_hd__xor2_2 _10436_ (.A(\term_mid[42] ),
    .B(\term_high[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01603_));
 sky130_fd_sc_hd__a22o_2 _10437_ (.A1(\term_mid[40] ),
    .A2(\term_high[40] ),
    .B1(\term_mid[41] ),
    .B2(\term_high[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01604_));
 sky130_fd_sc_hd__o21a_2 _10438_ (.A1(\term_mid[41] ),
    .A2(\term_high[41] ),
    .B1(_01604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01605_));
 sky130_fd_sc_hd__a31o_2 _10439_ (.A1(_01595_),
    .A2(_01599_),
    .A3(_01590_),
    .B1(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01606_));
 sky130_fd_sc_hd__a311o_2 _10440_ (.A1(_01595_),
    .A2(_01599_),
    .A3(_01590_),
    .B1(_01603_),
    .C1(_01605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01607_));
 sky130_fd_sc_hd__nand2_2 _10441_ (.A(_01606_),
    .B(_01603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01608_));
 sky130_fd_sc_hd__and3_2 _10442_ (.A(_09690_),
    .B(_01607_),
    .C(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00058_));
 sky130_fd_sc_hd__xor2_2 _10443_ (.A(\term_mid[43] ),
    .B(\term_high[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01609_));
 sky130_fd_sc_hd__a21bo_2 _10444_ (.A1(\term_mid[42] ),
    .A2(\term_high[42] ),
    .B1_N(_01608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01610_));
 sky130_fd_sc_hd__a21oi_2 _10445_ (.A1(_01610_),
    .A2(_01609_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01611_));
 sky130_fd_sc_hd__o21a_2 _10446_ (.A1(_01609_),
    .A2(_01610_),
    .B1(_01611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00059_));
 sky130_fd_sc_hd__xor2_2 _10447_ (.A(\term_mid[44] ),
    .B(\term_high[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01612_));
 sky130_fd_sc_hd__and3_2 _10448_ (.A(_01603_),
    .B(_01605_),
    .C(_01609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01613_));
 sky130_fd_sc_hd__o211a_2 _10449_ (.A1(\term_mid[43] ),
    .A2(\term_high[43] ),
    .B1(\term_mid[42] ),
    .C1(\term_high[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01614_));
 sky130_fd_sc_hd__a211o_2 _10450_ (.A1(\term_mid[43] ),
    .A2(\term_high[43] ),
    .B1(_01613_),
    .C1(_01614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01615_));
 sky130_fd_sc_hd__and4_2 _10451_ (.A(_01590_),
    .B(_01599_),
    .C(_01603_),
    .D(_01609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01616_));
 sky130_fd_sc_hd__a21o_2 _10452_ (.A1(_01595_),
    .A2(_01616_),
    .B1(_01615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01617_));
 sky130_fd_sc_hd__a211o_2 _10453_ (.A1(_01595_),
    .A2(_01616_),
    .B1(_01615_),
    .C1(_01612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01618_));
 sky130_fd_sc_hd__nand2_2 _10454_ (.A(_01617_),
    .B(_01612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01619_));
 sky130_fd_sc_hd__and3_2 _10455_ (.A(_09690_),
    .B(_01618_),
    .C(_01619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00060_));
 sky130_fd_sc_hd__xor2_2 _10456_ (.A(\term_mid[45] ),
    .B(\term_high[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01620_));
 sky130_fd_sc_hd__a21bo_2 _10457_ (.A1(\term_mid[44] ),
    .A2(\term_high[44] ),
    .B1_N(_01619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01621_));
 sky130_fd_sc_hd__a21oi_2 _10458_ (.A1(_01621_),
    .A2(_01620_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01622_));
 sky130_fd_sc_hd__o21a_2 _10459_ (.A1(_01620_),
    .A2(_01621_),
    .B1(_01622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_2 _10460_ (.A1(\term_mid[44] ),
    .A2(\term_high[44] ),
    .B1(\term_mid[45] ),
    .B2(\term_high[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01623_));
 sky130_fd_sc_hd__o21a_2 _10461_ (.A1(\term_mid[45] ),
    .A2(\term_high[45] ),
    .B1(_01623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01624_));
 sky130_fd_sc_hd__a31oi_2 _10462_ (.A1(_01617_),
    .A2(_01620_),
    .A3(_01612_),
    .B1(_01624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01625_));
 sky130_fd_sc_hd__and2_2 _10463_ (.A(\term_mid[46] ),
    .B(\term_high[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01626_));
 sky130_fd_sc_hd__nor2_2 _10464_ (.A(\term_mid[46] ),
    .B(\term_high[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_2 _10465_ (.A(_01626_),
    .B(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01628_));
 sky130_fd_sc_hd__o21a_2 _10466_ (.A1(_01626_),
    .A2(_01627_),
    .B1(_01625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01629_));
 sky130_fd_sc_hd__nor3_2 _10467_ (.A(_01625_),
    .B(_01626_),
    .C(_01627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01630_));
 sky130_fd_sc_hd__nor3_2 _10468_ (.A(rst),
    .B(_01629_),
    .C(_01630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00062_));
 sky130_fd_sc_hd__xor2_2 _10469_ (.A(\term_mid[47] ),
    .B(\term_high[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01631_));
 sky130_fd_sc_hd__a21o_2 _10470_ (.A1(\term_mid[46] ),
    .A2(\term_high[46] ),
    .B1(_01631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01632_));
 sky130_fd_sc_hd__o21ai_2 _10471_ (.A1(_01626_),
    .A2(_01630_),
    .B1(_01631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01633_));
 sky130_fd_sc_hd__o211a_2 _10472_ (.A1(_01632_),
    .A2(_01630_),
    .B1(_09690_),
    .C1(_01633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00063_));
 sky130_fd_sc_hd__nor2_2 _10473_ (.A(\term_mid[48] ),
    .B(\term_high[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01634_));
 sky130_fd_sc_hd__and2_2 _10474_ (.A(\term_mid[48] ),
    .B(\term_high[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01635_));
 sky130_fd_sc_hd__nor2_2 _10475_ (.A(_01634_),
    .B(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01636_));
 sky130_fd_sc_hd__and3_2 _10476_ (.A(_01624_),
    .B(_01628_),
    .C(_01631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01637_));
 sky130_fd_sc_hd__o211a_2 _10477_ (.A1(\term_mid[47] ),
    .A2(\term_high[47] ),
    .B1(\term_mid[46] ),
    .C1(\term_high[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01638_));
 sky130_fd_sc_hd__a211o_2 _10478_ (.A1(\term_mid[47] ),
    .A2(\term_high[47] ),
    .B1(_01637_),
    .C1(_01638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01639_));
 sky130_fd_sc_hd__a2111o_2 _10479_ (.A1(\term_mid[43] ),
    .A2(\term_high[43] ),
    .B1(_01613_),
    .C1(_01614_),
    .D1(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01640_));
 sky130_fd_sc_hd__a21o_2 _10480_ (.A1(_01595_),
    .A2(_01616_),
    .B1(_01640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01641_));
 sky130_fd_sc_hd__a41o_2 _10481_ (.A1(_01612_),
    .A2(_01620_),
    .A3(_01628_),
    .A4(_01631_),
    .B1(_01639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01642_));
 sky130_fd_sc_hd__a2bb2o_2 _10482_ (.A1_N(_01634_),
    .A2_N(_01635_),
    .B1(_01641_),
    .B2(_01642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01643_));
 sky130_fd_sc_hd__a31o_2 _10483_ (.A1(_01641_),
    .A2(_01642_),
    .A3(_01636_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01644_));
 sky130_fd_sc_hd__and2b_2 _10484_ (.A_N(_01644_),
    .B(_01643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00064_));
 sky130_fd_sc_hd__a31o_2 _10485_ (.A1(_01641_),
    .A2(_01642_),
    .A3(_01636_),
    .B1(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01645_));
 sky130_fd_sc_hd__a21oi_2 _10486_ (.A1(_01645_),
    .A2(\term_high[49] ),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01646_));
 sky130_fd_sc_hd__o21a_2 _10487_ (.A1(\term_high[49] ),
    .A2(_01645_),
    .B1(_01646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00065_));
 sky130_fd_sc_hd__a21oi_2 _10488_ (.A1(_01645_),
    .A2(\term_high[49] ),
    .B1(\term_high[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01647_));
 sky130_fd_sc_hd__a31o_2 _10489_ (.A1(_01645_),
    .A2(\term_high[50] ),
    .A3(\term_high[49] ),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01648_));
 sky130_fd_sc_hd__nor2_2 _10490_ (.A(_01647_),
    .B(_01648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00066_));
 sky130_fd_sc_hd__a31o_2 _10491_ (.A1(_01645_),
    .A2(\term_high[50] ),
    .A3(\term_high[49] ),
    .B1(\term_high[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01649_));
 sky130_fd_sc_hd__o2111a_2 _10492_ (.A1(\term_mid[48] ),
    .A2(\term_high[48] ),
    .B1(\term_high[49] ),
    .C1(\term_high[50] ),
    .D1(\term_high[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01650_));
 sky130_fd_sc_hd__nand3_2 _10493_ (.A(_01641_),
    .B(_01642_),
    .C(_01650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01651_));
 sky130_fd_sc_hd__nand4_2 _10494_ (.A(\term_high[49] ),
    .B(\term_high[50] ),
    .C(\term_high[51] ),
    .D(_01635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_2 _10495_ (.A(_01651_),
    .B(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01653_));
 sky130_fd_sc_hd__and4_2 _10496_ (.A(_09690_),
    .B(_01649_),
    .C(_01651_),
    .D(_01652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00067_));
 sky130_fd_sc_hd__a21oi_2 _10497_ (.A1(_01653_),
    .A2(\term_high[52] ),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01654_));
 sky130_fd_sc_hd__o21a_2 _10498_ (.A1(\term_high[52] ),
    .A2(_01653_),
    .B1(_01654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00068_));
 sky130_fd_sc_hd__a21oi_2 _10499_ (.A1(_01653_),
    .A2(\term_high[52] ),
    .B1(\term_high[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01655_));
 sky130_fd_sc_hd__and3_2 _10500_ (.A(_01653_),
    .B(\term_high[53] ),
    .C(\term_high[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01656_));
 sky130_fd_sc_hd__nor3_2 _10501_ (.A(rst),
    .B(_01655_),
    .C(_01656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00069_));
 sky130_fd_sc_hd__and3_2 _10502_ (.A(\term_high[52] ),
    .B(\term_high[53] ),
    .C(\term_high[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01657_));
 sky130_fd_sc_hd__a21oi_2 _10503_ (.A1(_01653_),
    .A2(_01657_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01658_));
 sky130_fd_sc_hd__o21a_2 _10504_ (.A1(\term_high[54] ),
    .A2(_01656_),
    .B1(_01658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00070_));
 sky130_fd_sc_hd__a21oi_2 _10505_ (.A1(_01653_),
    .A2(_01657_),
    .B1(\term_high[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01659_));
 sky130_fd_sc_hd__and3_2 _10506_ (.A(_01653_),
    .B(_01657_),
    .C(\term_high[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01660_));
 sky130_fd_sc_hd__nor3_2 _10507_ (.A(rst),
    .B(_01659_),
    .C(_01660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00071_));
 sky130_fd_sc_hd__a21oi_2 _10508_ (.A1(\term_high[56] ),
    .A2(_01660_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01661_));
 sky130_fd_sc_hd__o21a_2 _10509_ (.A1(\term_high[56] ),
    .A2(_01660_),
    .B1(_01661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00072_));
 sky130_fd_sc_hd__a21oi_2 _10510_ (.A1(\term_high[56] ),
    .A2(_01660_),
    .B1(\term_high[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01662_));
 sky130_fd_sc_hd__a311oi_2 _10511_ (.A1(\term_high[56] ),
    .A2(\term_high[57] ),
    .A3(_01660_),
    .B1(_01662_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00073_));
 sky130_fd_sc_hd__a31o_2 _10512_ (.A1(\term_high[56] ),
    .A2(\term_high[57] ),
    .A3(_01660_),
    .B1(\term_high[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01663_));
 sky130_fd_sc_hd__and3_2 _10513_ (.A(\term_high[56] ),
    .B(\term_high[57] ),
    .C(\term_high[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01664_));
 sky130_fd_sc_hd__nand4_2 _10514_ (.A(_01653_),
    .B(_01657_),
    .C(_01664_),
    .D(\term_high[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01665_));
 sky130_fd_sc_hd__and3_2 _10515_ (.A(_09690_),
    .B(_01663_),
    .C(_01665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00074_));
 sky130_fd_sc_hd__a21oi_2 _10516_ (.A1(_01660_),
    .A2(_01664_),
    .B1(\term_high[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01666_));
 sky130_fd_sc_hd__a311oi_2 _10517_ (.A1(\term_high[59] ),
    .A2(_01660_),
    .A3(_01664_),
    .B1(_01666_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00075_));
 sky130_fd_sc_hd__a31o_2 _10518_ (.A1(\term_high[59] ),
    .A2(_01660_),
    .A3(_01664_),
    .B1(\term_high[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01667_));
 sky130_fd_sc_hd__nand2_2 _10519_ (.A(\term_high[59] ),
    .B(\term_high[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_2 _10520_ (.A(_01665_),
    .B(_01668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01669_));
 sky130_fd_sc_hd__o211a_2 _10521_ (.A1(_01665_),
    .A2(_01668_),
    .B1(_01667_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00076_));
 sky130_fd_sc_hd__a21oi_2 _10522_ (.A1(\term_high[61] ),
    .A2(_01669_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01670_));
 sky130_fd_sc_hd__o21a_2 _10523_ (.A1(\term_high[61] ),
    .A2(_01669_),
    .B1(_01670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00077_));
 sky130_fd_sc_hd__a21oi_2 _10524_ (.A1(\term_high[61] ),
    .A2(_01669_),
    .B1(\term_high[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01671_));
 sky130_fd_sc_hd__a311oi_2 _10525_ (.A1(\term_high[61] ),
    .A2(\term_high[62] ),
    .A3(_01669_),
    .B1(_01671_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00078_));
 sky130_fd_sc_hd__a31oi_2 _10526_ (.A1(\term_high[61] ),
    .A2(\term_high[62] ),
    .A3(_01669_),
    .B1(\term_high[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01672_));
 sky130_fd_sc_hd__a41o_2 _10527_ (.A1(\term_high[61] ),
    .A2(\term_high[62] ),
    .A3(\term_high[63] ),
    .A4(_01669_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01673_));
 sky130_fd_sc_hd__nor2_2 _10528_ (.A(_01672_),
    .B(_01673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00079_));
 sky130_fd_sc_hd__and2_2 _10529_ (.A(_09690_),
    .B(\p_hh_pipe[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00080_));
 sky130_fd_sc_hd__and2_2 _10530_ (.A(_09690_),
    .B(\p_hh_pipe[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00081_));
 sky130_fd_sc_hd__and2_2 _10531_ (.A(_09690_),
    .B(\p_hh_pipe[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00082_));
 sky130_fd_sc_hd__and2_2 _10532_ (.A(_09690_),
    .B(\p_hh_pipe[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00083_));
 sky130_fd_sc_hd__and2_2 _10533_ (.A(_09690_),
    .B(\p_hh_pipe[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00084_));
 sky130_fd_sc_hd__and2_2 _10534_ (.A(_09690_),
    .B(\p_hh_pipe[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00085_));
 sky130_fd_sc_hd__and2_2 _10535_ (.A(_09690_),
    .B(\p_hh_pipe[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00086_));
 sky130_fd_sc_hd__and2_2 _10536_ (.A(_09690_),
    .B(\p_hh_pipe[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00087_));
 sky130_fd_sc_hd__and2_2 _10537_ (.A(_09690_),
    .B(\p_hh_pipe[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00088_));
 sky130_fd_sc_hd__and2_2 _10538_ (.A(_09690_),
    .B(\p_hh_pipe[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00089_));
 sky130_fd_sc_hd__and2_2 _10539_ (.A(_09690_),
    .B(\p_hh_pipe[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00090_));
 sky130_fd_sc_hd__and2_2 _10540_ (.A(_09690_),
    .B(\p_hh_pipe[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00091_));
 sky130_fd_sc_hd__and2_2 _10541_ (.A(_09690_),
    .B(\p_hh_pipe[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00092_));
 sky130_fd_sc_hd__and2_2 _10542_ (.A(_09690_),
    .B(\p_hh_pipe[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00093_));
 sky130_fd_sc_hd__and2_2 _10543_ (.A(_09690_),
    .B(\p_hh_pipe[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00094_));
 sky130_fd_sc_hd__and2_2 _10544_ (.A(_09690_),
    .B(\p_hh_pipe[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00095_));
 sky130_fd_sc_hd__and2_2 _10545_ (.A(_09690_),
    .B(\p_hh_pipe[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00096_));
 sky130_fd_sc_hd__and2_2 _10546_ (.A(_09690_),
    .B(\p_hh_pipe[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00097_));
 sky130_fd_sc_hd__and2_2 _10547_ (.A(_09690_),
    .B(\p_hh_pipe[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00098_));
 sky130_fd_sc_hd__and2_2 _10548_ (.A(_09690_),
    .B(\p_hh_pipe[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00099_));
 sky130_fd_sc_hd__and2_2 _10549_ (.A(_09690_),
    .B(\p_hh_pipe[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00100_));
 sky130_fd_sc_hd__and2_2 _10550_ (.A(_09690_),
    .B(\p_hh_pipe[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00101_));
 sky130_fd_sc_hd__and2_2 _10551_ (.A(_09690_),
    .B(\p_hh_pipe[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00102_));
 sky130_fd_sc_hd__and2_2 _10552_ (.A(_09690_),
    .B(\p_hh_pipe[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00103_));
 sky130_fd_sc_hd__and2_2 _10553_ (.A(_09690_),
    .B(\p_hh_pipe[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00104_));
 sky130_fd_sc_hd__and2_2 _10554_ (.A(_09690_),
    .B(\p_hh_pipe[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00105_));
 sky130_fd_sc_hd__and2_2 _10555_ (.A(_09690_),
    .B(\p_hh_pipe[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00106_));
 sky130_fd_sc_hd__and2_2 _10556_ (.A(_09690_),
    .B(\p_hh_pipe[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00107_));
 sky130_fd_sc_hd__and2_2 _10557_ (.A(_09690_),
    .B(\p_hh_pipe[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00108_));
 sky130_fd_sc_hd__and2_2 _10558_ (.A(_09690_),
    .B(\p_hh_pipe[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00109_));
 sky130_fd_sc_hd__and2_2 _10559_ (.A(_09690_),
    .B(\p_hh_pipe[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00110_));
 sky130_fd_sc_hd__and2_2 _10560_ (.A(_09690_),
    .B(\p_hh_pipe[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00111_));
 sky130_fd_sc_hd__and2_2 _10561_ (.A(_09690_),
    .B(\mid_sum[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00112_));
 sky130_fd_sc_hd__and2_2 _10562_ (.A(_09690_),
    .B(\mid_sum[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00113_));
 sky130_fd_sc_hd__and2_2 _10563_ (.A(_09690_),
    .B(\mid_sum[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00114_));
 sky130_fd_sc_hd__and2_2 _10564_ (.A(_09690_),
    .B(\mid_sum[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00115_));
 sky130_fd_sc_hd__and2_2 _10565_ (.A(_09690_),
    .B(\mid_sum[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00116_));
 sky130_fd_sc_hd__and2_2 _10566_ (.A(_09690_),
    .B(\mid_sum[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00117_));
 sky130_fd_sc_hd__and2_2 _10567_ (.A(_09690_),
    .B(\mid_sum[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00118_));
 sky130_fd_sc_hd__and2_2 _10568_ (.A(_09690_),
    .B(\mid_sum[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00119_));
 sky130_fd_sc_hd__and2_2 _10569_ (.A(_09690_),
    .B(\mid_sum[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00120_));
 sky130_fd_sc_hd__and2_2 _10570_ (.A(_09690_),
    .B(\mid_sum[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00121_));
 sky130_fd_sc_hd__and2_2 _10571_ (.A(_09690_),
    .B(\mid_sum[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00122_));
 sky130_fd_sc_hd__and2_2 _10572_ (.A(_09690_),
    .B(\mid_sum[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00123_));
 sky130_fd_sc_hd__and2_2 _10573_ (.A(_09690_),
    .B(\mid_sum[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00124_));
 sky130_fd_sc_hd__and2_2 _10574_ (.A(_09690_),
    .B(\mid_sum[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00125_));
 sky130_fd_sc_hd__and2_2 _10575_ (.A(_09690_),
    .B(\mid_sum[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00126_));
 sky130_fd_sc_hd__and2_2 _10576_ (.A(_09690_),
    .B(\mid_sum[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00127_));
 sky130_fd_sc_hd__and2_2 _10577_ (.A(_09690_),
    .B(\mid_sum[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00128_));
 sky130_fd_sc_hd__and2_2 _10578_ (.A(_09690_),
    .B(\mid_sum[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00129_));
 sky130_fd_sc_hd__and2_2 _10579_ (.A(_09690_),
    .B(\mid_sum[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00130_));
 sky130_fd_sc_hd__and2_2 _10580_ (.A(_09690_),
    .B(\mid_sum[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00131_));
 sky130_fd_sc_hd__and2_2 _10581_ (.A(_09690_),
    .B(\mid_sum[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00132_));
 sky130_fd_sc_hd__and2_2 _10582_ (.A(_09690_),
    .B(\mid_sum[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00133_));
 sky130_fd_sc_hd__and2_2 _10583_ (.A(_09690_),
    .B(\mid_sum[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00134_));
 sky130_fd_sc_hd__and2_2 _10584_ (.A(_09690_),
    .B(\mid_sum[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00135_));
 sky130_fd_sc_hd__and2_2 _10585_ (.A(_09690_),
    .B(\mid_sum[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00136_));
 sky130_fd_sc_hd__and2_2 _10586_ (.A(_09690_),
    .B(\mid_sum[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00137_));
 sky130_fd_sc_hd__and2_2 _10587_ (.A(_09690_),
    .B(\mid_sum[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00138_));
 sky130_fd_sc_hd__and2_2 _10588_ (.A(_09690_),
    .B(\mid_sum[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00139_));
 sky130_fd_sc_hd__and2_2 _10589_ (.A(_09690_),
    .B(\mid_sum[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00140_));
 sky130_fd_sc_hd__and2_2 _10590_ (.A(_09690_),
    .B(\mid_sum[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00141_));
 sky130_fd_sc_hd__and2_2 _10591_ (.A(_09690_),
    .B(\mid_sum[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00142_));
 sky130_fd_sc_hd__and2_2 _10592_ (.A(_09690_),
    .B(\mid_sum[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00143_));
 sky130_fd_sc_hd__and2_2 _10593_ (.A(_09690_),
    .B(\mid_sum[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00144_));
 sky130_fd_sc_hd__and2_2 _10594_ (.A(_09690_),
    .B(\p_ll_pipe[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00145_));
 sky130_fd_sc_hd__and2_2 _10595_ (.A(_09690_),
    .B(\p_ll_pipe[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00146_));
 sky130_fd_sc_hd__and2_2 _10596_ (.A(_09690_),
    .B(\p_ll_pipe[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00147_));
 sky130_fd_sc_hd__and2_2 _10597_ (.A(_09690_),
    .B(\p_ll_pipe[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00148_));
 sky130_fd_sc_hd__and2_2 _10598_ (.A(_09690_),
    .B(\p_ll_pipe[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00149_));
 sky130_fd_sc_hd__and2_2 _10599_ (.A(_09690_),
    .B(\p_ll_pipe[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00150_));
 sky130_fd_sc_hd__and2_2 _10600_ (.A(_09690_),
    .B(\p_ll_pipe[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00151_));
 sky130_fd_sc_hd__and2_2 _10601_ (.A(_09690_),
    .B(\p_ll_pipe[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00152_));
 sky130_fd_sc_hd__and2_2 _10602_ (.A(_09690_),
    .B(\p_ll_pipe[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00153_));
 sky130_fd_sc_hd__and2_2 _10603_ (.A(_09690_),
    .B(\p_ll_pipe[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00154_));
 sky130_fd_sc_hd__and2_2 _10604_ (.A(_09690_),
    .B(\p_ll_pipe[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00155_));
 sky130_fd_sc_hd__and2_2 _10605_ (.A(_09690_),
    .B(\p_ll_pipe[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00156_));
 sky130_fd_sc_hd__and2_2 _10606_ (.A(_09690_),
    .B(\p_ll_pipe[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00157_));
 sky130_fd_sc_hd__and2_2 _10607_ (.A(_09690_),
    .B(\p_ll_pipe[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00158_));
 sky130_fd_sc_hd__and2_2 _10608_ (.A(_09690_),
    .B(\p_ll_pipe[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00159_));
 sky130_fd_sc_hd__and2_2 _10609_ (.A(_09690_),
    .B(\p_ll_pipe[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00160_));
 sky130_fd_sc_hd__and2_2 _10610_ (.A(_09690_),
    .B(\p_ll_pipe[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00161_));
 sky130_fd_sc_hd__and2_2 _10611_ (.A(_09690_),
    .B(\p_ll_pipe[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00162_));
 sky130_fd_sc_hd__and2_2 _10612_ (.A(_09690_),
    .B(\p_ll_pipe[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00163_));
 sky130_fd_sc_hd__and2_2 _10613_ (.A(_09690_),
    .B(\p_ll_pipe[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00164_));
 sky130_fd_sc_hd__and2_2 _10614_ (.A(_09690_),
    .B(\p_ll_pipe[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00165_));
 sky130_fd_sc_hd__and2_2 _10615_ (.A(_09690_),
    .B(\p_ll_pipe[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00166_));
 sky130_fd_sc_hd__and2_2 _10616_ (.A(_09690_),
    .B(\p_ll_pipe[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00167_));
 sky130_fd_sc_hd__and2_2 _10617_ (.A(_09690_),
    .B(\p_ll_pipe[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00168_));
 sky130_fd_sc_hd__and2_2 _10618_ (.A(_09690_),
    .B(\p_ll_pipe[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00169_));
 sky130_fd_sc_hd__and2_2 _10619_ (.A(_09690_),
    .B(\p_ll_pipe[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00170_));
 sky130_fd_sc_hd__and2_2 _10620_ (.A(_09690_),
    .B(\p_ll_pipe[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00171_));
 sky130_fd_sc_hd__and2_2 _10621_ (.A(_09690_),
    .B(\p_ll_pipe[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00172_));
 sky130_fd_sc_hd__and2_2 _10622_ (.A(_09690_),
    .B(\p_ll_pipe[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00173_));
 sky130_fd_sc_hd__and2_2 _10623_ (.A(_09690_),
    .B(\p_ll_pipe[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00174_));
 sky130_fd_sc_hd__and2_2 _10624_ (.A(_09690_),
    .B(\p_ll_pipe[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00175_));
 sky130_fd_sc_hd__and2_2 _10625_ (.A(_09690_),
    .B(\p_ll_pipe[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00176_));
 sky130_fd_sc_hd__a21oi_2 _10626_ (.A1(\p_hl[0] ),
    .A2(\p_lh[0] ),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01674_));
 sky130_fd_sc_hd__o21a_2 _10627_ (.A1(\p_hl[0] ),
    .A2(\p_lh[0] ),
    .B1(_01674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00177_));
 sky130_fd_sc_hd__and2_2 _10628_ (.A(\p_hl[1] ),
    .B(\p_lh[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01675_));
 sky130_fd_sc_hd__nand2_2 _10629_ (.A(\p_hl[1] ),
    .B(\p_lh[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01676_));
 sky130_fd_sc_hd__nor2_2 _10630_ (.A(\p_hl[1] ),
    .B(\p_lh[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01677_));
 sky130_fd_sc_hd__o211ai_2 _10631_ (.A1(\p_hl[1] ),
    .A2(\p_lh[1] ),
    .B1(\p_hl[0] ),
    .C1(\p_lh[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01678_));
 sky130_fd_sc_hd__a2bb2o_2 _10632_ (.A1_N(_01675_),
    .A2_N(_01677_),
    .B1(\p_hl[0] ),
    .B2(\p_lh[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01679_));
 sky130_fd_sc_hd__o211a_2 _10633_ (.A1(_01678_),
    .A2(_01675_),
    .B1(_09690_),
    .C1(_01679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00178_));
 sky130_fd_sc_hd__nand2_2 _10634_ (.A(\p_hl[2] ),
    .B(\p_lh[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01680_));
 sky130_fd_sc_hd__and2b_2 _10635_ (.A_N(\p_hl[2] ),
    .B(\p_lh[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01681_));
 sky130_fd_sc_hd__and2b_2 _10636_ (.A_N(\p_lh[2] ),
    .B(\p_hl[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01682_));
 sky130_fd_sc_hd__nor2_2 _10637_ (.A(_01681_),
    .B(_01682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01683_));
 sky130_fd_sc_hd__o2bb2ai_2 _10638_ (.A1_N(_01676_),
    .A2_N(_01678_),
    .B1(_01681_),
    .B2(_01682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01684_));
 sky130_fd_sc_hd__a31o_2 _10639_ (.A1(_01676_),
    .A2(_01678_),
    .A3(_01683_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01685_));
 sky130_fd_sc_hd__and2b_2 _10640_ (.A_N(_01685_),
    .B(_01684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00179_));
 sky130_fd_sc_hd__nor2_2 _10641_ (.A(\p_hl[3] ),
    .B(\p_lh[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01686_));
 sky130_fd_sc_hd__and2_2 _10642_ (.A(\p_hl[3] ),
    .B(\p_lh[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01687_));
 sky130_fd_sc_hd__nor2_2 _10643_ (.A(_01686_),
    .B(_01687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01688_));
 sky130_fd_sc_hd__o211a_2 _10644_ (.A1(_01686_),
    .A2(_01687_),
    .B1(_01680_),
    .C1(_01684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01689_));
 sky130_fd_sc_hd__a21boi_2 _10645_ (.A1(_01680_),
    .A2(_01684_),
    .B1_N(_01688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01690_));
 sky130_fd_sc_hd__nor3_2 _10646_ (.A(rst),
    .B(_01689_),
    .C(_01690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00180_));
 sky130_fd_sc_hd__nor2_2 _10647_ (.A(\p_hl[4] ),
    .B(\p_lh[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01691_));
 sky130_fd_sc_hd__and2_2 _10648_ (.A(\p_hl[4] ),
    .B(\p_lh[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_2 _10649_ (.A(\p_hl[4] ),
    .B(\p_lh[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01693_));
 sky130_fd_sc_hd__a21oi_2 _10650_ (.A1(\p_hl[3] ),
    .A2(\p_lh[3] ),
    .B1(_01690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01694_));
 sky130_fd_sc_hd__o21ai_2 _10651_ (.A1(_01691_),
    .A2(_01692_),
    .B1(_01694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01695_));
 sky130_fd_sc_hd__or3_2 _10652_ (.A(_01691_),
    .B(_01692_),
    .C(_01694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01696_));
 sky130_fd_sc_hd__and3_2 _10653_ (.A(_09690_),
    .B(_01695_),
    .C(_01696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00181_));
 sky130_fd_sc_hd__o22ai_2 _10654_ (.A1(\p_hl[4] ),
    .A2(\p_lh[4] ),
    .B1(_01687_),
    .B2(_01690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01697_));
 sky130_fd_sc_hd__o21ai_2 _10655_ (.A1(_01691_),
    .A2(_01694_),
    .B1(_01693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_2 _10656_ (.A(\p_hl[5] ),
    .B(\p_lh[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01699_));
 sky130_fd_sc_hd__or2_2 _10657_ (.A(\p_hl[5] ),
    .B(\p_lh[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01700_));
 sky130_fd_sc_hd__a21oi_2 _10658_ (.A1(_01699_),
    .A2(_01700_),
    .B1(_01698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01701_));
 sky130_fd_sc_hd__a31o_2 _10659_ (.A1(_01698_),
    .A2(_01699_),
    .A3(_01700_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01702_));
 sky130_fd_sc_hd__nor2_2 _10660_ (.A(_01701_),
    .B(_01702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00182_));
 sky130_fd_sc_hd__nor2_2 _10661_ (.A(_09537_),
    .B(_09548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01703_));
 sky130_fd_sc_hd__nor2_2 _10662_ (.A(\p_hl[6] ),
    .B(\p_lh[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01704_));
 sky130_fd_sc_hd__nand3_2 _10663_ (.A(_01693_),
    .B(_01697_),
    .C(_01699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01705_));
 sky130_fd_sc_hd__o21ai_2 _10664_ (.A1(\p_hl[5] ),
    .A2(\p_lh[5] ),
    .B1(_01705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01706_));
 sky130_fd_sc_hd__a2bb2o_2 _10665_ (.A1_N(_01703_),
    .A2_N(_01704_),
    .B1(_01705_),
    .B2(_01700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01707_));
 sky130_fd_sc_hd__or3_2 _10666_ (.A(_01703_),
    .B(_01704_),
    .C(_01706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01708_));
 sky130_fd_sc_hd__and3_2 _10667_ (.A(_09690_),
    .B(_01707_),
    .C(_01708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_2 _10668_ (.A(\p_hl[7] ),
    .B(\p_lh[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01709_));
 sky130_fd_sc_hd__or2_2 _10669_ (.A(\p_hl[7] ),
    .B(\p_lh[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01710_));
 sky130_fd_sc_hd__o211ai_2 _10670_ (.A1(\p_hl[6] ),
    .A2(\p_lh[6] ),
    .B1(_01700_),
    .C1(_01705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01711_));
 sky130_fd_sc_hd__o21ai_2 _10671_ (.A1(_09537_),
    .A2(_09548_),
    .B1(_01711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01712_));
 sky130_fd_sc_hd__a21oi_2 _10672_ (.A1(_01709_),
    .A2(_01710_),
    .B1(_01712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01713_));
 sky130_fd_sc_hd__a31o_2 _10673_ (.A1(_01712_),
    .A2(_01710_),
    .A3(_01709_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01714_));
 sky130_fd_sc_hd__nor2_2 _10674_ (.A(_01713_),
    .B(_01714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00184_));
 sky130_fd_sc_hd__o211ai_2 _10675_ (.A1(_09537_),
    .A2(_09548_),
    .B1(_01709_),
    .C1(_01711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_2 _10676_ (.A(\p_hl[8] ),
    .B(\p_lh[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01716_));
 sky130_fd_sc_hd__xor2_2 _10677_ (.A(\p_hl[8] ),
    .B(\p_lh[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01717_));
 sky130_fd_sc_hd__a21oi_2 _10678_ (.A1(_01710_),
    .A2(_01715_),
    .B1(_01717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01718_));
 sky130_fd_sc_hd__o211ai_2 _10679_ (.A1(\p_hl[7] ),
    .A2(\p_lh[7] ),
    .B1(_01717_),
    .C1(_01715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01719_));
 sky130_fd_sc_hd__a311oi_2 _10680_ (.A1(_01710_),
    .A2(_01717_),
    .A3(_01715_),
    .B1(rst),
    .C1(_01718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00185_));
 sky130_fd_sc_hd__xnor2_2 _10681_ (.A(\p_hl[9] ),
    .B(\p_lh[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01720_));
 sky130_fd_sc_hd__a21oi_2 _10682_ (.A1(_01716_),
    .A2(_01719_),
    .B1(_01720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01721_));
 sky130_fd_sc_hd__a31o_2 _10683_ (.A1(_01716_),
    .A2(_01719_),
    .A3(_01720_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01722_));
 sky130_fd_sc_hd__nor2_2 _10684_ (.A(_01721_),
    .B(_01722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00186_));
 sky130_fd_sc_hd__nor2_2 _10685_ (.A(\p_hl[10] ),
    .B(\p_lh[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_2 _10686_ (.A(\p_hl[10] ),
    .B(\p_lh[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01724_));
 sky130_fd_sc_hd__and2b_2 _10687_ (.A_N(_01723_),
    .B(_01724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01725_));
 sky130_fd_sc_hd__o211ai_2 _10688_ (.A1(_09559_),
    .A2(_09570_),
    .B1(_01716_),
    .C1(_01719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01726_));
 sky130_fd_sc_hd__o21a_2 _10689_ (.A1(\p_hl[9] ),
    .A2(\p_lh[9] ),
    .B1(_01726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01727_));
 sky130_fd_sc_hd__o211ai_2 _10690_ (.A1(\p_hl[9] ),
    .A2(\p_lh[9] ),
    .B1(_01725_),
    .C1(_01726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01728_));
 sky130_fd_sc_hd__o21ai_2 _10691_ (.A1(_01725_),
    .A2(_01727_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01729_));
 sky130_fd_sc_hd__a21oi_2 _10692_ (.A1(_01725_),
    .A2(_01727_),
    .B1(_01729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00187_));
 sky130_fd_sc_hd__nor2_2 _10693_ (.A(\p_hl[11] ),
    .B(\p_lh[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01730_));
 sky130_fd_sc_hd__and2_2 _10694_ (.A(\p_hl[11] ),
    .B(\p_lh[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_2 _10695_ (.A(\p_hl[11] ),
    .B(\p_lh[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01732_));
 sky130_fd_sc_hd__o211ai_2 _10696_ (.A1(_01730_),
    .A2(_01731_),
    .B1(_01724_),
    .C1(_01728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01733_));
 sky130_fd_sc_hd__a211o_2 _10697_ (.A1(_01724_),
    .A2(_01728_),
    .B1(_01730_),
    .C1(_01731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01734_));
 sky130_fd_sc_hd__and3_2 _10698_ (.A(_09690_),
    .B(_01733_),
    .C(_01734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00188_));
 sky130_fd_sc_hd__nor2_2 _10699_ (.A(\p_hl[12] ),
    .B(\p_lh[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01735_));
 sky130_fd_sc_hd__and2_2 _10700_ (.A(\p_hl[12] ),
    .B(\p_lh[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01736_));
 sky130_fd_sc_hd__nor2_2 _10701_ (.A(_01735_),
    .B(_01736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01737_));
 sky130_fd_sc_hd__nand3_2 _10702_ (.A(_01724_),
    .B(_01728_),
    .C(_01732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01738_));
 sky130_fd_sc_hd__o21a_2 _10703_ (.A1(\p_hl[11] ),
    .A2(\p_lh[11] ),
    .B1(_01738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01739_));
 sky130_fd_sc_hd__o211ai_2 _10704_ (.A1(\p_hl[11] ),
    .A2(\p_lh[11] ),
    .B1(_01737_),
    .C1(_01738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01740_));
 sky130_fd_sc_hd__a21oi_2 _10705_ (.A1(_01739_),
    .A2(_01737_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01741_));
 sky130_fd_sc_hd__o21a_2 _10706_ (.A1(_01737_),
    .A2(_01739_),
    .B1(_01741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00189_));
 sky130_fd_sc_hd__a21o_2 _10707_ (.A1(_01739_),
    .A2(_01737_),
    .B1(_01736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01742_));
 sky130_fd_sc_hd__nand2_2 _10708_ (.A(\p_hl[13] ),
    .B(\p_lh[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01743_));
 sky130_fd_sc_hd__or2_2 _10709_ (.A(\p_hl[13] ),
    .B(\p_lh[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01744_));
 sky130_fd_sc_hd__a21oi_2 _10710_ (.A1(_01743_),
    .A2(_01744_),
    .B1(_01742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01745_));
 sky130_fd_sc_hd__a31o_2 _10711_ (.A1(_01742_),
    .A2(_01743_),
    .A3(_01744_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01746_));
 sky130_fd_sc_hd__nor2_2 _10712_ (.A(_01745_),
    .B(_01746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00190_));
 sky130_fd_sc_hd__xor2_2 _10713_ (.A(\p_hl[14] ),
    .B(\p_lh[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01747_));
 sky130_fd_sc_hd__nand3b_2 _10714_ (.A_N(_01736_),
    .B(_01740_),
    .C(_01743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01748_));
 sky130_fd_sc_hd__o21a_2 _10715_ (.A1(\p_hl[13] ),
    .A2(\p_lh[13] ),
    .B1(_01748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01749_));
 sky130_fd_sc_hd__a31o_2 _10716_ (.A1(_01744_),
    .A2(_01748_),
    .A3(_01747_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01750_));
 sky130_fd_sc_hd__o21ba_2 _10717_ (.A1(_01747_),
    .A2(_01749_),
    .B1_N(_01750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00191_));
 sky130_fd_sc_hd__xor2_2 _10718_ (.A(\p_hl[15] ),
    .B(\p_lh[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01751_));
 sky130_fd_sc_hd__a32o_2 _10719_ (.A1(_01744_),
    .A2(_01748_),
    .A3(_01747_),
    .B1(\p_hl[14] ),
    .B2(\p_lh[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01752_));
 sky130_fd_sc_hd__a21oi_2 _10720_ (.A1(_01752_),
    .A2(_01751_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01753_));
 sky130_fd_sc_hd__o21a_2 _10721_ (.A1(_01751_),
    .A2(_01752_),
    .B1(_01753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00192_));
 sky130_fd_sc_hd__xnor2_2 _10722_ (.A(\p_hl[16] ),
    .B(\p_lh[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01754_));
 sky130_fd_sc_hd__and2_2 _10723_ (.A(_01747_),
    .B(_01751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01755_));
 sky130_fd_sc_hd__o211ai_2 _10724_ (.A1(\p_hl[13] ),
    .A2(\p_lh[13] ),
    .B1(_01755_),
    .C1(_01748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01756_));
 sky130_fd_sc_hd__o211a_2 _10725_ (.A1(\p_hl[15] ),
    .A2(\p_lh[15] ),
    .B1(\p_hl[14] ),
    .C1(\p_lh[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01757_));
 sky130_fd_sc_hd__a21oi_2 _10726_ (.A1(\p_hl[15] ),
    .A2(\p_lh[15] ),
    .B1(_01757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_2 _10727_ (.A(_01756_),
    .B(_01758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01759_));
 sky130_fd_sc_hd__a21oi_2 _10728_ (.A1(_01756_),
    .A2(_01758_),
    .B1(_01754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01760_));
 sky130_fd_sc_hd__a31o_2 _10729_ (.A1(_01754_),
    .A2(_01756_),
    .A3(_01758_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01761_));
 sky130_fd_sc_hd__nor2_2 _10730_ (.A(_01760_),
    .B(_01761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00193_));
 sky130_fd_sc_hd__xor2_2 _10731_ (.A(\p_hl[17] ),
    .B(\p_lh[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01762_));
 sky130_fd_sc_hd__a21o_2 _10732_ (.A1(\p_hl[16] ),
    .A2(\p_lh[16] ),
    .B1(_01760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01763_));
 sky130_fd_sc_hd__a21oi_2 _10733_ (.A1(_01763_),
    .A2(_01762_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01764_));
 sky130_fd_sc_hd__o21a_2 _10734_ (.A1(_01762_),
    .A2(_01763_),
    .B1(_01764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00194_));
 sky130_fd_sc_hd__nor2_2 _10735_ (.A(\p_hl[18] ),
    .B(\p_lh[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01765_));
 sky130_fd_sc_hd__and2_2 _10736_ (.A(\p_hl[18] ),
    .B(\p_lh[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01766_));
 sky130_fd_sc_hd__nor2_2 _10737_ (.A(_01765_),
    .B(_01766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01767_));
 sky130_fd_sc_hd__nand3b_2 _10738_ (.A_N(_01754_),
    .B(_01759_),
    .C(_01762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01768_));
 sky130_fd_sc_hd__a22o_2 _10739_ (.A1(\p_hl[16] ),
    .A2(\p_lh[16] ),
    .B1(\p_hl[17] ),
    .B2(\p_lh[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01769_));
 sky130_fd_sc_hd__o21ai_2 _10740_ (.A1(\p_hl[17] ),
    .A2(\p_lh[17] ),
    .B1(_01769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01770_));
 sky130_fd_sc_hd__nand2_2 _10741_ (.A(_01768_),
    .B(_01770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01771_));
 sky130_fd_sc_hd__a211oi_2 _10742_ (.A1(_01768_),
    .A2(_01770_),
    .B1(_01765_),
    .C1(_01766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01772_));
 sky130_fd_sc_hd__a21oi_2 _10743_ (.A1(_01771_),
    .A2(_01767_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01773_));
 sky130_fd_sc_hd__o21a_2 _10744_ (.A1(_01767_),
    .A2(_01771_),
    .B1(_01773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00195_));
 sky130_fd_sc_hd__xor2_2 _10745_ (.A(\p_hl[19] ),
    .B(\p_lh[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01774_));
 sky130_fd_sc_hd__or3_2 _10746_ (.A(_01766_),
    .B(_01772_),
    .C(_01774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01775_));
 sky130_fd_sc_hd__o21ai_2 _10747_ (.A1(_01766_),
    .A2(_01772_),
    .B1(_01774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01776_));
 sky130_fd_sc_hd__and3_2 _10748_ (.A(_09690_),
    .B(_01775_),
    .C(_01776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00196_));
 sky130_fd_sc_hd__nor2_2 _10749_ (.A(\p_hl[20] ),
    .B(\p_lh[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01777_));
 sky130_fd_sc_hd__and2_2 _10750_ (.A(\p_hl[20] ),
    .B(\p_lh[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01778_));
 sky130_fd_sc_hd__nor2_2 _10751_ (.A(_01777_),
    .B(_01778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01779_));
 sky130_fd_sc_hd__o211a_2 _10752_ (.A1(\p_hl[19] ),
    .A2(\p_lh[19] ),
    .B1(\p_hl[18] ),
    .C1(\p_lh[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01780_));
 sky130_fd_sc_hd__o211a_2 _10753_ (.A1(\p_hl[17] ),
    .A2(\p_lh[17] ),
    .B1(_01769_),
    .C1(_01774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01781_));
 sky130_fd_sc_hd__a221o_2 _10754_ (.A1(\p_hl[19] ),
    .A2(\p_lh[19] ),
    .B1(_01767_),
    .B2(_01781_),
    .C1(_01780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01782_));
 sky130_fd_sc_hd__and4b_2 _10755_ (.A_N(_01754_),
    .B(_01762_),
    .C(_01767_),
    .D(_01774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01783_));
 sky130_fd_sc_hd__a21boi_2 _10756_ (.A1(_01756_),
    .A2(_01758_),
    .B1_N(_01783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01784_));
 sky130_fd_sc_hd__a21o_2 _10757_ (.A1(_01759_),
    .A2(_01783_),
    .B1(_01782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01785_));
 sky130_fd_sc_hd__a21oi_2 _10758_ (.A1(_01759_),
    .A2(_01783_),
    .B1(_01782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01786_));
 sky130_fd_sc_hd__o21a_2 _10759_ (.A1(_01782_),
    .A2(_01784_),
    .B1(_01779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01787_));
 sky130_fd_sc_hd__o31a_2 _10760_ (.A1(_01777_),
    .A2(_01778_),
    .A3(_01786_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01788_));
 sky130_fd_sc_hd__o31a_2 _10761_ (.A1(_01779_),
    .A2(_01782_),
    .A3(_01784_),
    .B1(_01788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00197_));
 sky130_fd_sc_hd__xor2_2 _10762_ (.A(\p_hl[21] ),
    .B(\p_lh[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01789_));
 sky130_fd_sc_hd__a221o_2 _10763_ (.A1(\p_hl[20] ),
    .A2(\p_lh[20] ),
    .B1(_01779_),
    .B2(_01785_),
    .C1(_01789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01790_));
 sky130_fd_sc_hd__o21ai_2 _10764_ (.A1(_01778_),
    .A2(_01787_),
    .B1(_01789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01791_));
 sky130_fd_sc_hd__and3_2 _10765_ (.A(_09690_),
    .B(_01790_),
    .C(_01791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00198_));
 sky130_fd_sc_hd__and2_2 _10766_ (.A(\p_hl[22] ),
    .B(\p_lh[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01792_));
 sky130_fd_sc_hd__nor2_2 _10767_ (.A(\p_hl[22] ),
    .B(\p_lh[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_2 _10768_ (.A(_01792_),
    .B(_01793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01794_));
 sky130_fd_sc_hd__a22o_2 _10769_ (.A1(\p_hl[20] ),
    .A2(\p_lh[20] ),
    .B1(\p_hl[21] ),
    .B2(\p_lh[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01795_));
 sky130_fd_sc_hd__o21a_2 _10770_ (.A1(\p_hl[21] ),
    .A2(\p_lh[21] ),
    .B1(_01795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01796_));
 sky130_fd_sc_hd__a21oi_2 _10771_ (.A1(_01787_),
    .A2(_01789_),
    .B1(_01796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01797_));
 sky130_fd_sc_hd__a31o_2 _10772_ (.A1(_01779_),
    .A2(_01785_),
    .A3(_01789_),
    .B1(_01796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01798_));
 sky130_fd_sc_hd__nor3_2 _10773_ (.A(_01792_),
    .B(_01793_),
    .C(_01797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01799_));
 sky130_fd_sc_hd__o31a_2 _10774_ (.A1(_01792_),
    .A2(_01793_),
    .A3(_01797_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01800_));
 sky130_fd_sc_hd__o21a_2 _10775_ (.A1(_01794_),
    .A2(_01798_),
    .B1(_01800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00199_));
 sky130_fd_sc_hd__nor2_2 _10776_ (.A(\p_hl[23] ),
    .B(\p_lh[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01801_));
 sky130_fd_sc_hd__and2_2 _10777_ (.A(\p_hl[23] ),
    .B(\p_lh[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01802_));
 sky130_fd_sc_hd__nor2_2 _10778_ (.A(_01801_),
    .B(_01802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01803_));
 sky130_fd_sc_hd__or3_2 _10779_ (.A(_01792_),
    .B(_01799_),
    .C(_01803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01804_));
 sky130_fd_sc_hd__o21ai_2 _10780_ (.A1(_01792_),
    .A2(_01799_),
    .B1(_01803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01805_));
 sky130_fd_sc_hd__and3_2 _10781_ (.A(_09690_),
    .B(_01804_),
    .C(_01805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00200_));
 sky130_fd_sc_hd__and2_2 _10782_ (.A(\p_hl[24] ),
    .B(\p_lh[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_2 _10783_ (.A(\p_hl[24] ),
    .B(\p_lh[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01807_));
 sky130_fd_sc_hd__or2_2 _10784_ (.A(_01806_),
    .B(_01807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01808_));
 sky130_fd_sc_hd__o211a_2 _10785_ (.A1(\p_hl[23] ),
    .A2(\p_lh[23] ),
    .B1(\p_hl[22] ),
    .C1(\p_lh[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01809_));
 sky130_fd_sc_hd__nand4_2 _10786_ (.A(_01779_),
    .B(_01789_),
    .C(_01794_),
    .D(_01803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01810_));
 sky130_fd_sc_hd__o21bai_2 _10787_ (.A1(_01782_),
    .A2(_01784_),
    .B1_N(_01810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01811_));
 sky130_fd_sc_hd__a311oi_2 _10788_ (.A1(_01794_),
    .A2(_01796_),
    .A3(_01803_),
    .B1(_01809_),
    .C1(_01802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_2 _10789_ (.A(_01811_),
    .B(_01812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01813_));
 sky130_fd_sc_hd__o21a_2 _10790_ (.A1(_01786_),
    .A2(_01810_),
    .B1(_01812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01814_));
 sky130_fd_sc_hd__a21oi_2 _10791_ (.A1(_01808_),
    .A2(_01814_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01815_));
 sky130_fd_sc_hd__o31a_2 _10792_ (.A1(_01806_),
    .A2(_01807_),
    .A3(_01814_),
    .B1(_01815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00201_));
 sky130_fd_sc_hd__nor2_2 _10793_ (.A(\p_hl[25] ),
    .B(\p_lh[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01816_));
 sky130_fd_sc_hd__and2_2 _10794_ (.A(\p_hl[25] ),
    .B(\p_lh[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01817_));
 sky130_fd_sc_hd__nor2_2 _10795_ (.A(_01816_),
    .B(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01818_));
 sky130_fd_sc_hd__o21bai_2 _10796_ (.A1(_01808_),
    .A2(_01814_),
    .B1_N(_01806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01819_));
 sky130_fd_sc_hd__a21oi_2 _10797_ (.A1(_01819_),
    .A2(_01818_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01820_));
 sky130_fd_sc_hd__o21a_2 _10798_ (.A1(_01818_),
    .A2(_01819_),
    .B1(_01820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00202_));
 sky130_fd_sc_hd__xor2_2 _10799_ (.A(\p_hl[26] ),
    .B(\p_lh[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01821_));
 sky130_fd_sc_hd__a21oi_2 _10800_ (.A1(\p_hl[25] ),
    .A2(\p_lh[25] ),
    .B1(_01806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01822_));
 sky130_fd_sc_hd__or4_2 _10801_ (.A(_01806_),
    .B(_01807_),
    .C(_01816_),
    .D(_01817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01823_));
 sky130_fd_sc_hd__o22ai_2 _10802_ (.A1(_01816_),
    .A2(_01822_),
    .B1(_01823_),
    .B2(_01814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01824_));
 sky130_fd_sc_hd__or2_2 _10803_ (.A(_01821_),
    .B(_01824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01825_));
 sky130_fd_sc_hd__nand2_2 _10804_ (.A(_01824_),
    .B(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01826_));
 sky130_fd_sc_hd__and3_2 _10805_ (.A(_09690_),
    .B(_01825_),
    .C(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00203_));
 sky130_fd_sc_hd__xor2_2 _10806_ (.A(\p_hl[27] ),
    .B(\p_lh[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01827_));
 sky130_fd_sc_hd__a21bo_2 _10807_ (.A1(\p_hl[26] ),
    .A2(\p_lh[26] ),
    .B1_N(_01826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01828_));
 sky130_fd_sc_hd__a21oi_2 _10808_ (.A1(_01828_),
    .A2(_01827_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01829_));
 sky130_fd_sc_hd__o21a_2 _10809_ (.A1(_01827_),
    .A2(_01828_),
    .B1(_01829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00204_));
 sky130_fd_sc_hd__nor2_2 _10810_ (.A(\p_hl[28] ),
    .B(\p_lh[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01830_));
 sky130_fd_sc_hd__and2_2 _10811_ (.A(\p_hl[28] ),
    .B(\p_lh[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01831_));
 sky130_fd_sc_hd__nor2_2 _10812_ (.A(_01830_),
    .B(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01832_));
 sky130_fd_sc_hd__and4b_2 _10813_ (.A_N(_01808_),
    .B(_01818_),
    .C(_01821_),
    .D(_01827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01833_));
 sky130_fd_sc_hd__and4bb_2 _10814_ (.A_N(_01816_),
    .B_N(_01822_),
    .C(_01827_),
    .D(_01821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01834_));
 sky130_fd_sc_hd__o211a_2 _10815_ (.A1(\p_hl[27] ),
    .A2(\p_lh[27] ),
    .B1(\p_hl[26] ),
    .C1(\p_lh[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01835_));
 sky130_fd_sc_hd__a211o_2 _10816_ (.A1(\p_hl[27] ),
    .A2(\p_lh[27] ),
    .B1(_01834_),
    .C1(_01835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01836_));
 sky130_fd_sc_hd__a21o_2 _10817_ (.A1(_01813_),
    .A2(_01833_),
    .B1(_01836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01837_));
 sky130_fd_sc_hd__a21oi_2 _10818_ (.A1(_01837_),
    .A2(_01832_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01838_));
 sky130_fd_sc_hd__o21a_2 _10819_ (.A1(_01832_),
    .A2(_01837_),
    .B1(_01838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00205_));
 sky130_fd_sc_hd__xor2_2 _10820_ (.A(\p_hl[29] ),
    .B(\p_lh[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01839_));
 sky130_fd_sc_hd__a21o_2 _10821_ (.A1(_01837_),
    .A2(_01832_),
    .B1(_01831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01840_));
 sky130_fd_sc_hd__o21ai_2 _10822_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01841_));
 sky130_fd_sc_hd__a21oi_2 _10823_ (.A1(_01839_),
    .A2(_01840_),
    .B1(_01841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00206_));
 sky130_fd_sc_hd__xnor2_2 _10824_ (.A(\p_hl[30] ),
    .B(\p_lh[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01842_));
 sky130_fd_sc_hd__and2_2 _10825_ (.A(_01832_),
    .B(_01839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01843_));
 sky130_fd_sc_hd__o211a_2 _10826_ (.A1(\p_hl[29] ),
    .A2(\p_lh[29] ),
    .B1(\p_hl[28] ),
    .C1(\p_lh[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01844_));
 sky130_fd_sc_hd__a21o_2 _10827_ (.A1(\p_hl[29] ),
    .A2(\p_lh[29] ),
    .B1(_01844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01845_));
 sky130_fd_sc_hd__a21oi_2 _10828_ (.A1(_01837_),
    .A2(_01843_),
    .B1(_01845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_2 _10829_ (.A(_01842_),
    .B(_01846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01847_));
 sky130_fd_sc_hd__o21ai_2 _10830_ (.A1(_01842_),
    .A2(_01846_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01848_));
 sky130_fd_sc_hd__a21oi_2 _10831_ (.A1(_01842_),
    .A2(_01846_),
    .B1(_01848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00207_));
 sky130_fd_sc_hd__nor2_2 _10832_ (.A(\p_hl[31] ),
    .B(\p_lh[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01849_));
 sky130_fd_sc_hd__and2_2 _10833_ (.A(\p_hl[31] ),
    .B(\p_lh[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01850_));
 sky130_fd_sc_hd__or2_2 _10834_ (.A(_01849_),
    .B(_01850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01851_));
 sky130_fd_sc_hd__a21oi_2 _10835_ (.A1(\p_hl[30] ),
    .A2(\p_lh[30] ),
    .B1(_01847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01852_));
 sky130_fd_sc_hd__a2bb2o_2 _10836_ (.A1_N(_01849_),
    .A2_N(_01850_),
    .B1(\p_hl[30] ),
    .B2(\p_lh[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01853_));
 sky130_fd_sc_hd__o221a_2 _10837_ (.A1(_01847_),
    .A2(_01853_),
    .B1(_01851_),
    .B2(_01852_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_2 _10838_ (.A1(\p_hl[30] ),
    .A2(\p_lh[30] ),
    .B1(\p_hl[31] ),
    .B2(\p_lh[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01854_));
 sky130_fd_sc_hd__o221a_2 _10839_ (.A1(\p_hl[31] ),
    .A2(\p_lh[31] ),
    .B1(_01854_),
    .B2(_01847_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00209_));
 sky130_fd_sc_hd__and2_2 _10840_ (.A(_09690_),
    .B(\p_hh[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00210_));
 sky130_fd_sc_hd__and2_2 _10841_ (.A(_09690_),
    .B(\p_hh[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00211_));
 sky130_fd_sc_hd__and2_2 _10842_ (.A(_09690_),
    .B(\p_hh[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00212_));
 sky130_fd_sc_hd__and2_2 _10843_ (.A(_09690_),
    .B(\p_hh[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00213_));
 sky130_fd_sc_hd__and2_2 _10844_ (.A(_09690_),
    .B(\p_hh[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00214_));
 sky130_fd_sc_hd__and2_2 _10845_ (.A(_09690_),
    .B(\p_hh[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00215_));
 sky130_fd_sc_hd__and2_2 _10846_ (.A(_09690_),
    .B(\p_hh[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00216_));
 sky130_fd_sc_hd__and2_2 _10847_ (.A(_09690_),
    .B(\p_hh[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00217_));
 sky130_fd_sc_hd__and2_2 _10848_ (.A(_09690_),
    .B(\p_hh[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00218_));
 sky130_fd_sc_hd__and2_2 _10849_ (.A(_09690_),
    .B(\p_hh[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00219_));
 sky130_fd_sc_hd__and2_2 _10850_ (.A(_09690_),
    .B(\p_hh[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00220_));
 sky130_fd_sc_hd__and2_2 _10851_ (.A(_09690_),
    .B(\p_hh[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00221_));
 sky130_fd_sc_hd__and2_2 _10852_ (.A(_09690_),
    .B(\p_hh[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00222_));
 sky130_fd_sc_hd__and2_2 _10853_ (.A(_09690_),
    .B(\p_hh[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00223_));
 sky130_fd_sc_hd__and2_2 _10854_ (.A(_09690_),
    .B(\p_hh[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00224_));
 sky130_fd_sc_hd__and2_2 _10855_ (.A(_09690_),
    .B(\p_hh[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00225_));
 sky130_fd_sc_hd__and2_2 _10856_ (.A(_09690_),
    .B(\p_hh[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00226_));
 sky130_fd_sc_hd__and2_2 _10857_ (.A(_09690_),
    .B(\p_hh[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00227_));
 sky130_fd_sc_hd__and2_2 _10858_ (.A(_09690_),
    .B(\p_hh[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00228_));
 sky130_fd_sc_hd__and2_2 _10859_ (.A(_09690_),
    .B(\p_hh[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00229_));
 sky130_fd_sc_hd__and2_2 _10860_ (.A(_09690_),
    .B(\p_hh[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00230_));
 sky130_fd_sc_hd__and2_2 _10861_ (.A(_09690_),
    .B(\p_hh[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00231_));
 sky130_fd_sc_hd__and2_2 _10862_ (.A(_09690_),
    .B(\p_hh[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00232_));
 sky130_fd_sc_hd__and2_2 _10863_ (.A(_09690_),
    .B(\p_hh[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00233_));
 sky130_fd_sc_hd__and2_2 _10864_ (.A(_09690_),
    .B(\p_hh[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00234_));
 sky130_fd_sc_hd__and2_2 _10865_ (.A(_09690_),
    .B(\p_hh[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00235_));
 sky130_fd_sc_hd__and2_2 _10866_ (.A(_09690_),
    .B(\p_hh[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00236_));
 sky130_fd_sc_hd__and2_2 _10867_ (.A(_09690_),
    .B(\p_hh[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00237_));
 sky130_fd_sc_hd__and2_2 _10868_ (.A(_09690_),
    .B(\p_hh[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00238_));
 sky130_fd_sc_hd__and2_2 _10869_ (.A(_09690_),
    .B(\p_hh[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00239_));
 sky130_fd_sc_hd__and2_2 _10870_ (.A(_09690_),
    .B(\p_hh[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00240_));
 sky130_fd_sc_hd__and2_2 _10871_ (.A(_09690_),
    .B(\p_hh[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00241_));
 sky130_fd_sc_hd__and2_2 _10872_ (.A(_09690_),
    .B(\p_ll[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00242_));
 sky130_fd_sc_hd__and2_2 _10873_ (.A(_09690_),
    .B(\p_ll[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00243_));
 sky130_fd_sc_hd__and2_2 _10874_ (.A(_09690_),
    .B(\p_ll[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00244_));
 sky130_fd_sc_hd__and2_2 _10875_ (.A(_09690_),
    .B(\p_ll[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00245_));
 sky130_fd_sc_hd__and2_2 _10876_ (.A(_09690_),
    .B(\p_ll[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00246_));
 sky130_fd_sc_hd__and2_2 _10877_ (.A(_09690_),
    .B(\p_ll[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00247_));
 sky130_fd_sc_hd__and2_2 _10878_ (.A(_09690_),
    .B(\p_ll[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00248_));
 sky130_fd_sc_hd__and2_2 _10879_ (.A(_09690_),
    .B(\p_ll[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00249_));
 sky130_fd_sc_hd__and2_2 _10880_ (.A(_09690_),
    .B(\p_ll[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00250_));
 sky130_fd_sc_hd__and2_2 _10881_ (.A(_09690_),
    .B(\p_ll[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00251_));
 sky130_fd_sc_hd__and2_2 _10882_ (.A(_09690_),
    .B(\p_ll[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00252_));
 sky130_fd_sc_hd__and2_2 _10883_ (.A(_09690_),
    .B(\p_ll[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00253_));
 sky130_fd_sc_hd__and2_2 _10884_ (.A(_09690_),
    .B(\p_ll[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00254_));
 sky130_fd_sc_hd__and2_2 _10885_ (.A(_09690_),
    .B(\p_ll[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00255_));
 sky130_fd_sc_hd__and2_2 _10886_ (.A(_09690_),
    .B(\p_ll[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00256_));
 sky130_fd_sc_hd__and2_2 _10887_ (.A(_09690_),
    .B(\p_ll[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00257_));
 sky130_fd_sc_hd__and2_2 _10888_ (.A(_09690_),
    .B(\p_ll[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00258_));
 sky130_fd_sc_hd__and2_2 _10889_ (.A(_09690_),
    .B(\p_ll[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00259_));
 sky130_fd_sc_hd__and2_2 _10890_ (.A(_09690_),
    .B(\p_ll[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00260_));
 sky130_fd_sc_hd__and2_2 _10891_ (.A(_09690_),
    .B(\p_ll[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00261_));
 sky130_fd_sc_hd__and2_2 _10892_ (.A(_09690_),
    .B(\p_ll[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00262_));
 sky130_fd_sc_hd__and2_2 _10893_ (.A(_09690_),
    .B(\p_ll[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00263_));
 sky130_fd_sc_hd__and2_2 _10894_ (.A(_09690_),
    .B(\p_ll[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00264_));
 sky130_fd_sc_hd__and2_2 _10895_ (.A(_09690_),
    .B(\p_ll[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00265_));
 sky130_fd_sc_hd__and2_2 _10896_ (.A(_09690_),
    .B(\p_ll[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00266_));
 sky130_fd_sc_hd__and2_2 _10897_ (.A(_09690_),
    .B(\p_ll[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00267_));
 sky130_fd_sc_hd__and2_2 _10898_ (.A(_09690_),
    .B(\p_ll[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00268_));
 sky130_fd_sc_hd__and2_2 _10899_ (.A(_09690_),
    .B(\p_ll[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00269_));
 sky130_fd_sc_hd__and2_2 _10900_ (.A(_09690_),
    .B(\p_ll[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00270_));
 sky130_fd_sc_hd__and2_2 _10901_ (.A(_09690_),
    .B(\p_ll[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00271_));
 sky130_fd_sc_hd__and2_2 _10902_ (.A(_09690_),
    .B(\p_ll[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00272_));
 sky130_fd_sc_hd__and2_2 _10903_ (.A(_09690_),
    .B(\p_ll[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00273_));
 sky130_fd_sc_hd__and3_2 _10904_ (.A(_09690_),
    .B(\b_h[0] ),
    .C(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00274_));
 sky130_fd_sc_hd__nand2_2 _10905_ (.A(\a_h[0] ),
    .B(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_2 _10906_ (.A(_09526_),
    .B(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_2 _10907_ (.A(\b_h[0] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01857_));
 sky130_fd_sc_hd__a22o_2 _10908_ (.A1(\a_h[1] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01858_));
 sky130_fd_sc_hd__o311a_2 _10909_ (.A1(_09526_),
    .A2(_09581_),
    .A3(_01855_),
    .B1(_01858_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00275_));
 sky130_fd_sc_hd__nand2_2 _10910_ (.A(\a_h[0] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_2 _10911_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01860_));
 sky130_fd_sc_hd__a22oi_2 _10912_ (.A1(\a_h[2] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01861_));
 sky130_fd_sc_hd__a31oi_2 _10913_ (.A1(\a_h[1] ),
    .A2(\a_h[2] ),
    .A3(_01856_),
    .B1(_01861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01862_));
 sky130_fd_sc_hd__xnor2_2 _10914_ (.A(_01859_),
    .B(_01862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01863_));
 sky130_fd_sc_hd__a31oi_2 _10915_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_01856_),
    .B1(_01863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01864_));
 sky130_fd_sc_hd__and4_2 _10916_ (.A(_01863_),
    .B(_01856_),
    .C(\a_h[1] ),
    .D(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01865_));
 sky130_fd_sc_hd__nor3_2 _10917_ (.A(rst),
    .B(_01864_),
    .C(_01865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00276_));
 sky130_fd_sc_hd__and2_2 _10918_ (.A(\a_h[0] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01866_));
 sky130_fd_sc_hd__o22ai_2 _10919_ (.A1(_01857_),
    .A2(_01860_),
    .B1(_01859_),
    .B2(_01861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_2 _10920_ (.A(\a_h[1] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01868_));
 sky130_fd_sc_hd__a22oi_2 _10921_ (.A1(\a_h[3] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01869_));
 sky130_fd_sc_hd__a22o_2 _10922_ (.A1(\a_h[3] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01870_));
 sky130_fd_sc_hd__nand2_2 _10923_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01871_));
 sky130_fd_sc_hd__nand4_2 _10924_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01872_));
 sky130_fd_sc_hd__a21o_2 _10925_ (.A1(_01870_),
    .A2(_01872_),
    .B1(_01868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01873_));
 sky130_fd_sc_hd__nand3_2 _10926_ (.A(_01868_),
    .B(_01870_),
    .C(_01872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01874_));
 sky130_fd_sc_hd__a21bo_2 _10927_ (.A1(_01873_),
    .A2(_01874_),
    .B1_N(_01867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01875_));
 sky130_fd_sc_hd__nand3b_2 _10928_ (.A_N(_01867_),
    .B(_01873_),
    .C(_01874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01876_));
 sky130_fd_sc_hd__a21oi_2 _10929_ (.A1(_01875_),
    .A2(_01876_),
    .B1(_01866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01877_));
 sky130_fd_sc_hd__and3_2 _10930_ (.A(_01876_),
    .B(\b_h[3] ),
    .C(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01878_));
 sky130_fd_sc_hd__nand2_2 _10931_ (.A(_01876_),
    .B(_01866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01879_));
 sky130_fd_sc_hd__a21oi_2 _10932_ (.A1(_01878_),
    .A2(_01875_),
    .B1(_01877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01880_));
 sky130_fd_sc_hd__a41o_2 _10933_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_01856_),
    .A4(_01863_),
    .B1(_01880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01881_));
 sky130_fd_sc_hd__nand2_2 _10934_ (.A(_01865_),
    .B(_01880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01882_));
 sky130_fd_sc_hd__and3_2 _10935_ (.A(_09690_),
    .B(_01881_),
    .C(_01882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00277_));
 sky130_fd_sc_hd__and3_2 _10936_ (.A(\a_h[1] ),
    .B(\b_h[4] ),
    .C(_01866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01883_));
 sky130_fd_sc_hd__a22oi_2 _10937_ (.A1(\a_h[1] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_2 _10938_ (.A(\a_h[2] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_2 _10939_ (.A(\a_h[3] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_2 _10940_ (.A(\a_h[4] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_2 _10941_ (.A(\a_h[3] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01888_));
 sky130_fd_sc_hd__nand4_2 _10942_ (.A(\a_h[3] ),
    .B(\a_h[4] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01889_));
 sky130_fd_sc_hd__a22oi_2 _10943_ (.A1(\a_h[4] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_2 _10944_ (.A(_01886_),
    .B(_01887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01891_));
 sky130_fd_sc_hd__a22o_2 _10945_ (.A1(\a_h[2] ),
    .A2(\b_h[2] ),
    .B1(_01889_),
    .B2(_01891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01892_));
 sky130_fd_sc_hd__nand4_2 _10946_ (.A(_01891_),
    .B(\b_h[2] ),
    .C(\a_h[2] ),
    .D(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01893_));
 sky130_fd_sc_hd__o21ai_2 _10947_ (.A1(_01868_),
    .A2(_01869_),
    .B1(_01872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01894_));
 sky130_fd_sc_hd__a21oi_2 _10948_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_01894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01895_));
 sky130_fd_sc_hd__a21o_2 _10949_ (.A1(_01892_),
    .A2(_01893_),
    .B1(_01894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01896_));
 sky130_fd_sc_hd__nand3_2 _10950_ (.A(_01892_),
    .B(_01893_),
    .C(_01894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01897_));
 sky130_fd_sc_hd__a211o_2 _10951_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_01883_),
    .C1(_01884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01898_));
 sky130_fd_sc_hd__o211ai_2 _10952_ (.A1(_01883_),
    .A2(_01884_),
    .B1(_01896_),
    .C1(_01897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01899_));
 sky130_fd_sc_hd__nand4_2 _10953_ (.A(_01875_),
    .B(_01879_),
    .C(_01898_),
    .D(_01899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01900_));
 sky130_fd_sc_hd__a22o_2 _10954_ (.A1(_01875_),
    .A2(_01879_),
    .B1(_01898_),
    .B2(_01899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01901_));
 sky130_fd_sc_hd__nand2_2 _10955_ (.A(_01900_),
    .B(_01901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01902_));
 sky130_fd_sc_hd__or2_2 _10956_ (.A(_01882_),
    .B(_01902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01903_));
 sky130_fd_sc_hd__a41o_2 _10957_ (.A1(_01901_),
    .A2(_01865_),
    .A3(_01900_),
    .A4(_01880_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01904_));
 sky130_fd_sc_hd__a21oi_2 _10958_ (.A1(_01882_),
    .A2(_01902_),
    .B1(_01904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00278_));
 sky130_fd_sc_hd__o21a_2 _10959_ (.A1(_01883_),
    .A2(_01884_),
    .B1(_01897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01905_));
 sky130_fd_sc_hd__nor2_2 _10960_ (.A(_01895_),
    .B(_01905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01906_));
 sky130_fd_sc_hd__nand2_2 _10961_ (.A(\a_h[0] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01907_));
 sky130_fd_sc_hd__a22oi_2 _10962_ (.A1(\a_h[2] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_2 _10963_ (.A(\a_h[2] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01909_));
 sky130_fd_sc_hd__and4_2 _10964_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01910_));
 sky130_fd_sc_hd__nand4_2 _10965_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01911_));
 sky130_fd_sc_hd__o21ai_2 _10966_ (.A1(_09177_),
    .A2(_09602_),
    .B1(_01911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01912_));
 sky130_fd_sc_hd__o21bai_2 _10967_ (.A1(_01908_),
    .A2(_01910_),
    .B1_N(_01907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01913_));
 sky130_fd_sc_hd__o21ai_2 _10968_ (.A1(_01908_),
    .A2(_01912_),
    .B1(_01913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01914_));
 sky130_fd_sc_hd__o21ai_2 _10969_ (.A1(_01885_),
    .A2(_01890_),
    .B1(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01915_));
 sky130_fd_sc_hd__o21a_2 _10970_ (.A1(_01885_),
    .A2(_01890_),
    .B1(_01889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01916_));
 sky130_fd_sc_hd__nand2_2 _10971_ (.A(\a_h[3] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_2 _10972_ (.A(\a_h[4] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_2 _10973_ (.A(\a_h[5] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01919_));
 sky130_fd_sc_hd__nand2_2 _10974_ (.A(_01918_),
    .B(_01919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01920_));
 sky130_fd_sc_hd__nand2_2 _10975_ (.A(\a_h[5] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01921_));
 sky130_fd_sc_hd__nand4_2 _10976_ (.A(\a_h[4] ),
    .B(\a_h[5] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01922_));
 sky130_fd_sc_hd__a22o_2 _10977_ (.A1(\a_h[3] ),
    .A2(\b_h[2] ),
    .B1(_01920_),
    .B2(_01922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01923_));
 sky130_fd_sc_hd__o2111ai_2 _10978_ (.A1(_01887_),
    .A2(_01921_),
    .B1(\a_h[3] ),
    .C1(\b_h[2] ),
    .D1(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01924_));
 sky130_fd_sc_hd__o221ai_2 _10979_ (.A1(_09406_),
    .A2(_09592_),
    .B1(_01887_),
    .B2(_01921_),
    .C1(_01920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01925_));
 sky130_fd_sc_hd__a21o_2 _10980_ (.A1(_01920_),
    .A2(_01922_),
    .B1(_01917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01926_));
 sky130_fd_sc_hd__nand3_2 _10981_ (.A(_01916_),
    .B(_01925_),
    .C(_01926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01927_));
 sky130_fd_sc_hd__nand3_2 _10982_ (.A(_01923_),
    .B(_01924_),
    .C(_01915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01928_));
 sky130_fd_sc_hd__o2111ai_2 _10983_ (.A1(_01908_),
    .A2(_01912_),
    .B1(_01913_),
    .C1(_01927_),
    .D1(_01928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01929_));
 sky130_fd_sc_hd__a21bo_2 _10984_ (.A1(_01927_),
    .A2(_01928_),
    .B1_N(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01930_));
 sky130_fd_sc_hd__nand3_2 _10985_ (.A(_01927_),
    .B(_01928_),
    .C(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01931_));
 sky130_fd_sc_hd__a21o_2 _10986_ (.A1(_01927_),
    .A2(_01928_),
    .B1(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01932_));
 sky130_fd_sc_hd__nand3_2 _10987_ (.A(_01906_),
    .B(_01931_),
    .C(_01932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01933_));
 sky130_fd_sc_hd__o211ai_2 _10988_ (.A1(_01895_),
    .A2(_01905_),
    .B1(_01929_),
    .C1(_01930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01934_));
 sky130_fd_sc_hd__a21boi_2 _10989_ (.A1(_01933_),
    .A2(_01934_),
    .B1_N(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01935_));
 sky130_fd_sc_hd__a31oi_2 _10990_ (.A1(_01932_),
    .A2(_01906_),
    .A3(_01931_),
    .B1(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01936_));
 sky130_fd_sc_hd__a31o_2 _10991_ (.A1(_01906_),
    .A2(_01931_),
    .A3(_01932_),
    .B1(_01883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01937_));
 sky130_fd_sc_hd__a21oi_2 _10992_ (.A1(_01934_),
    .A2(_01936_),
    .B1(_01935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01938_));
 sky130_fd_sc_hd__o211ai_2 _10993_ (.A1(_01882_),
    .A2(_01902_),
    .B1(_01938_),
    .C1(_01901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01939_));
 sky130_fd_sc_hd__or2_2 _10994_ (.A(_01901_),
    .B(_01938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01940_));
 sky130_fd_sc_hd__o2111a_2 _10995_ (.A1(_01938_),
    .A2(_01903_),
    .B1(_09690_),
    .C1(_01940_),
    .D1(_01939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00279_));
 sky130_fd_sc_hd__nand2_2 _10996_ (.A(_01927_),
    .B(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01941_));
 sky130_fd_sc_hd__a32oi_2 _10997_ (.A1(_01915_),
    .A2(_01923_),
    .A3(_01924_),
    .B1(_01927_),
    .B2(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01942_));
 sky130_fd_sc_hd__a32o_2 _10998_ (.A1(_01915_),
    .A2(_01923_),
    .A3(_01924_),
    .B1(_01927_),
    .B2(_01914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_2 _10999_ (.A(\a_h[1] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_2 _11000_ (.A(\a_h[3] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01945_));
 sky130_fd_sc_hd__nand2_2 _11001_ (.A(\a_h[3] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01946_));
 sky130_fd_sc_hd__nand4_2 _11002_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01947_));
 sky130_fd_sc_hd__a22oi_2 _11003_ (.A1(\a_h[3] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01948_));
 sky130_fd_sc_hd__nand2_2 _11004_ (.A(_01909_),
    .B(_01946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01949_));
 sky130_fd_sc_hd__nand3_2 _11005_ (.A(_01944_),
    .B(_01947_),
    .C(_01949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01950_));
 sky130_fd_sc_hd__a21o_2 _11006_ (.A1(_01947_),
    .A2(_01949_),
    .B1(_01944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01951_));
 sky130_fd_sc_hd__a22o_2 _11007_ (.A1(\a_h[1] ),
    .A2(\b_h[5] ),
    .B1(_01947_),
    .B2(_01949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01952_));
 sky130_fd_sc_hd__nand4_2 _11008_ (.A(_01949_),
    .B(\b_h[5] ),
    .C(\a_h[1] ),
    .D(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01953_));
 sky130_fd_sc_hd__nand2_2 _11009_ (.A(_01952_),
    .B(_01953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_2 _11010_ (.A(_01950_),
    .B(_01951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01955_));
 sky130_fd_sc_hd__a22o_2 _11011_ (.A1(_01918_),
    .A2(_01919_),
    .B1(_01922_),
    .B2(_01917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01956_));
 sky130_fd_sc_hd__a22oi_2 _11012_ (.A1(_01918_),
    .A2(_01919_),
    .B1(_01922_),
    .B2(_01917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01957_));
 sky130_fd_sc_hd__and2_2 _11013_ (.A(\a_h[4] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01958_));
 sky130_fd_sc_hd__nand2_2 _11014_ (.A(\a_h[4] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_2 _11015_ (.A(\a_h[6] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01960_));
 sky130_fd_sc_hd__nand2_2 _11016_ (.A(_01921_),
    .B(_01960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_2 _11017_ (.A(\a_h[6] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01962_));
 sky130_fd_sc_hd__nand4_2 _11018_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01963_));
 sky130_fd_sc_hd__a21oi_2 _11019_ (.A1(_01961_),
    .A2(_01963_),
    .B1(_01958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01964_));
 sky130_fd_sc_hd__a22o_2 _11020_ (.A1(\a_h[4] ),
    .A2(\b_h[2] ),
    .B1(_01961_),
    .B2(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01965_));
 sky130_fd_sc_hd__nand3_2 _11021_ (.A(_01961_),
    .B(_01963_),
    .C(_01958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01966_));
 sky130_fd_sc_hd__o221ai_2 _11022_ (.A1(_09417_),
    .A2(_09592_),
    .B1(_01919_),
    .B2(_01962_),
    .C1(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01967_));
 sky130_fd_sc_hd__a21o_2 _11023_ (.A1(_01961_),
    .A2(_01963_),
    .B1(_01959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01968_));
 sky130_fd_sc_hd__nand2_2 _11024_ (.A(_01957_),
    .B(_01966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_2 _11025_ (.A(_01964_),
    .B(_01969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01970_));
 sky130_fd_sc_hd__a21oi_2 _11026_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01971_));
 sky130_fd_sc_hd__nand3_2 _11027_ (.A(_01968_),
    .B(_01956_),
    .C(_01967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01972_));
 sky130_fd_sc_hd__o21ai_2 _11028_ (.A1(_01964_),
    .A2(_01969_),
    .B1(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01973_));
 sky130_fd_sc_hd__o2111ai_2 _11029_ (.A1(_01964_),
    .A2(_01969_),
    .B1(_01972_),
    .C1(_01953_),
    .D1(_01952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01974_));
 sky130_fd_sc_hd__o2bb2a_2 _11030_ (.A1_N(_01952_),
    .A2_N(_01953_),
    .B1(_01970_),
    .B2(_01971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01975_));
 sky130_fd_sc_hd__o21ai_2 _11031_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01976_));
 sky130_fd_sc_hd__nand2_2 _11032_ (.A(_01954_),
    .B(_01972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01977_));
 sky130_fd_sc_hd__o21ai_2 _11033_ (.A1(_01970_),
    .A2(_01971_),
    .B1(_01955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01978_));
 sky130_fd_sc_hd__o211ai_2 _11034_ (.A1(_01970_),
    .A2(_01977_),
    .B1(_01942_),
    .C1(_01978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01979_));
 sky130_fd_sc_hd__o2bb2ai_2 _11035_ (.A1_N(_01928_),
    .A2_N(_01941_),
    .B1(_01954_),
    .B2(_01973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01980_));
 sky130_fd_sc_hd__nand3_2 _11036_ (.A(_01943_),
    .B(_01974_),
    .C(_01976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01981_));
 sky130_fd_sc_hd__nand2_2 _11037_ (.A(\a_h[0] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01982_));
 sky130_fd_sc_hd__a21o_2 _11038_ (.A1(_01907_),
    .A2(_01911_),
    .B1(_01908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01983_));
 sky130_fd_sc_hd__and4b_2 _11039_ (.A_N(_01908_),
    .B(_01912_),
    .C(\a_h[0] ),
    .D(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01984_));
 sky130_fd_sc_hd__and2_2 _11040_ (.A(_01982_),
    .B(_01983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_2 _11041_ (.A(_01984_),
    .B(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01986_));
 sky130_fd_sc_hd__o211ai_2 _11042_ (.A1(_01980_),
    .A2(_01975_),
    .B1(_01979_),
    .C1(_01986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01987_));
 sky130_fd_sc_hd__o2bb2ai_2 _11043_ (.A1_N(_01979_),
    .A2_N(_01981_),
    .B1(_01984_),
    .B2(_01985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01988_));
 sky130_fd_sc_hd__a22oi_2 _11044_ (.A1(_01934_),
    .A2(_01937_),
    .B1(_01987_),
    .B2(_01988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01989_));
 sky130_fd_sc_hd__nor3_2 _11045_ (.A(_01901_),
    .B(_01938_),
    .C(_01989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01990_));
 sky130_fd_sc_hd__and4_2 _11046_ (.A(_01934_),
    .B(_01937_),
    .C(_01987_),
    .D(_01988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01991_));
 sky130_fd_sc_hd__nand4_2 _11047_ (.A(_01934_),
    .B(_01937_),
    .C(_01987_),
    .D(_01988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01992_));
 sky130_fd_sc_hd__nor4_2 _11048_ (.A(_01882_),
    .B(_01938_),
    .C(_01989_),
    .D(_01902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01993_));
 sky130_fd_sc_hd__a21o_2 _11049_ (.A1(_01993_),
    .A2(_01992_),
    .B1(_01990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01994_));
 sky130_fd_sc_hd__o221a_2 _11050_ (.A1(_01989_),
    .A2(_01991_),
    .B1(_01938_),
    .B2(_01903_),
    .C1(_01940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01995_));
 sky130_fd_sc_hd__nor3_2 _11051_ (.A(rst),
    .B(_01994_),
    .C(_01995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00280_));
 sky130_fd_sc_hd__o2bb2ai_2 _11052_ (.A1_N(_01986_),
    .A2_N(_01979_),
    .B1(_01975_),
    .B2(_01980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01996_));
 sky130_fd_sc_hd__a2bb2oi_2 _11053_ (.A1_N(_01975_),
    .A2_N(_01980_),
    .B1(_01986_),
    .B2(_01979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01997_));
 sky130_fd_sc_hd__a32oi_2 _11054_ (.A1(_01968_),
    .A2(_01956_),
    .A3(_01967_),
    .B1(_01951_),
    .B2(_01950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01998_));
 sky130_fd_sc_hd__a21oi_2 _11055_ (.A1(_01955_),
    .A2(_01972_),
    .B1(_01970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_2 _11056_ (.A(_01959_),
    .B(_01963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02000_));
 sky130_fd_sc_hd__nand2_2 _11057_ (.A(_01961_),
    .B(_02000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02001_));
 sky130_fd_sc_hd__a21boi_2 _11058_ (.A1(_01959_),
    .A2(_01963_),
    .B1_N(_01961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02002_));
 sky130_fd_sc_hd__nand2_2 _11059_ (.A(\a_h[5] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_2 _11060_ (.A(\a_h[7] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02004_));
 sky130_fd_sc_hd__a22o_2 _11061_ (.A1(\a_h[7] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02005_));
 sky130_fd_sc_hd__nand2_2 _11062_ (.A(\a_h[7] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02006_));
 sky130_fd_sc_hd__nand2_2 _11063_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02007_));
 sky130_fd_sc_hd__nand4_2 _11064_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02008_));
 sky130_fd_sc_hd__o2bb2ai_2 _11065_ (.A1_N(_01962_),
    .A2_N(_02004_),
    .B1(_02007_),
    .B2(_01857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02009_));
 sky130_fd_sc_hd__o21ai_2 _11066_ (.A1(_09428_),
    .A2(_09592_),
    .B1(_02009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02010_));
 sky130_fd_sc_hd__and4_2 _11067_ (.A(_02005_),
    .B(_02008_),
    .C(\a_h[5] ),
    .D(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02011_));
 sky130_fd_sc_hd__o2111ai_2 _11068_ (.A1(_01857_),
    .A2(_02007_),
    .B1(\a_h[5] ),
    .C1(\b_h[2] ),
    .D1(_02005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02012_));
 sky130_fd_sc_hd__o221ai_2 _11069_ (.A1(_09428_),
    .A2(_09592_),
    .B1(_01857_),
    .B2(_02007_),
    .C1(_02005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02013_));
 sky130_fd_sc_hd__nand3_2 _11070_ (.A(_02009_),
    .B(\b_h[2] ),
    .C(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02014_));
 sky130_fd_sc_hd__nand3_2 _11071_ (.A(_02014_),
    .B(_02001_),
    .C(_02013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02015_));
 sky130_fd_sc_hd__a21o_2 _11072_ (.A1(_02003_),
    .A2(_02009_),
    .B1(_02001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02016_));
 sky130_fd_sc_hd__nand3_2 _11073_ (.A(_02002_),
    .B(_02010_),
    .C(_02012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02017_));
 sky130_fd_sc_hd__and2_2 _11074_ (.A(\a_h[2] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02018_));
 sky130_fd_sc_hd__nand2_2 _11075_ (.A(\a_h[2] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_2 _11076_ (.A(\a_h[4] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02020_));
 sky130_fd_sc_hd__a22oi_2 _11077_ (.A1(\a_h[4] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_2 _11078_ (.A(_01945_),
    .B(_02020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02022_));
 sky130_fd_sc_hd__nand4_2 _11079_ (.A(\a_h[3] ),
    .B(\a_h[4] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02023_));
 sky130_fd_sc_hd__a21oi_2 _11080_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_02018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02024_));
 sky130_fd_sc_hd__and3_2 _11081_ (.A(_02022_),
    .B(_02023_),
    .C(_02018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02025_));
 sky130_fd_sc_hd__and3_2 _11082_ (.A(_02019_),
    .B(_02022_),
    .C(_02023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02026_));
 sky130_fd_sc_hd__a21oi_2 _11083_ (.A1(_02022_),
    .A2(_02023_),
    .B1(_02019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_2 _11084_ (.A(_02024_),
    .B(_02025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02028_));
 sky130_fd_sc_hd__o2bb2ai_2 _11085_ (.A1_N(_02015_),
    .A2_N(_02017_),
    .B1(_02026_),
    .B2(_02027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02029_));
 sky130_fd_sc_hd__o211ai_2 _11086_ (.A1(_02024_),
    .A2(_02025_),
    .B1(_02015_),
    .C1(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02030_));
 sky130_fd_sc_hd__o211ai_2 _11087_ (.A1(_02026_),
    .A2(_02027_),
    .B1(_02015_),
    .C1(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02031_));
 sky130_fd_sc_hd__o2bb2ai_2 _11088_ (.A1_N(_02015_),
    .A2_N(_02017_),
    .B1(_02024_),
    .B2(_02025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02032_));
 sky130_fd_sc_hd__a21oi_2 _11089_ (.A1(_02029_),
    .A2(_02030_),
    .B1(_01999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02033_));
 sky130_fd_sc_hd__o211ai_2 _11090_ (.A1(_01970_),
    .A2(_01998_),
    .B1(_02031_),
    .C1(_02032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02034_));
 sky130_fd_sc_hd__nand3_2 _11091_ (.A(_01999_),
    .B(_02029_),
    .C(_02030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02035_));
 sky130_fd_sc_hd__nand2_2 _11092_ (.A(_02034_),
    .B(_02035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_2 _11093_ (.A(\a_h[1] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02037_));
 sky130_fd_sc_hd__and4_2 _11094_ (.A(\a_h[0] ),
    .B(\a_h[1] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02038_));
 sky130_fd_sc_hd__a22oi_2 _11095_ (.A1(\a_h[1] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02039_));
 sky130_fd_sc_hd__or2_2 _11096_ (.A(_02038_),
    .B(_02039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02040_));
 sky130_fd_sc_hd__o21a_2 _11097_ (.A1(_01944_),
    .A2(_01948_),
    .B1(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02041_));
 sky130_fd_sc_hd__nor2_2 _11098_ (.A(_02040_),
    .B(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02042_));
 sky130_fd_sc_hd__inv_2 _11099_ (.A(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02043_));
 sky130_fd_sc_hd__o221a_2 _11100_ (.A1(_01948_),
    .A2(_01944_),
    .B1(_02039_),
    .B2(_02038_),
    .C1(_01947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02044_));
 sky130_fd_sc_hd__nor2_2 _11101_ (.A(_02042_),
    .B(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_2 _11102_ (.A(_02036_),
    .B(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02046_));
 sky130_fd_sc_hd__o211ai_2 _11103_ (.A1(_02042_),
    .A2(_02044_),
    .B1(_02034_),
    .C1(_02035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02047_));
 sky130_fd_sc_hd__o2bb2ai_2 _11104_ (.A1_N(_02034_),
    .A2_N(_02035_),
    .B1(_02042_),
    .B2(_02044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02048_));
 sky130_fd_sc_hd__inv_2 _11105_ (.A(_02048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02049_));
 sky130_fd_sc_hd__nand3_2 _11106_ (.A(_02034_),
    .B(_02035_),
    .C(_02045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_2 _11107_ (.A(_01996_),
    .B(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02051_));
 sky130_fd_sc_hd__nand3_2 _11108_ (.A(_01996_),
    .B(_02048_),
    .C(_02050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02052_));
 sky130_fd_sc_hd__nand3_2 _11109_ (.A(_01997_),
    .B(_02046_),
    .C(_02047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_2 _11110_ (.A(_02053_),
    .B(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02054_));
 sky130_fd_sc_hd__o211a_2 _11111_ (.A1(_01982_),
    .A2(_01983_),
    .B1(_02052_),
    .C1(_02053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02055_));
 sky130_fd_sc_hd__a21boi_2 _11112_ (.A1(_02052_),
    .A2(_02053_),
    .B1_N(_01984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_2 _11113_ (.A(_02055_),
    .B(_02056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02057_));
 sky130_fd_sc_hd__nor2_2 _11114_ (.A(_01991_),
    .B(_01994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02058_));
 sky130_fd_sc_hd__o41a_2 _11115_ (.A1(_01991_),
    .A2(_02055_),
    .A3(_02056_),
    .A4(_01994_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02059_));
 sky130_fd_sc_hd__o21ai_2 _11116_ (.A1(_02055_),
    .A2(_02056_),
    .B1(_01991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02060_));
 sky130_fd_sc_hd__o21a_2 _11117_ (.A1(_02057_),
    .A2(_02058_),
    .B1(_02059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00281_));
 sky130_fd_sc_hd__o2bb2ai_2 _11118_ (.A1_N(_02028_),
    .A2_N(_02015_),
    .B1(_02011_),
    .B2(_02016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02061_));
 sky130_fd_sc_hd__a21boi_2 _11119_ (.A1(_02028_),
    .A2(_02015_),
    .B1_N(_02017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_2 _11120_ (.A(\a_h[3] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02063_));
 sky130_fd_sc_hd__nand2_2 _11121_ (.A(\a_h[5] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02064_));
 sky130_fd_sc_hd__a22oi_2 _11122_ (.A1(\a_h[5] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02065_));
 sky130_fd_sc_hd__a22o_2 _11123_ (.A1(\a_h[5] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02066_));
 sky130_fd_sc_hd__nand2_2 _11124_ (.A(\a_h[5] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02067_));
 sky130_fd_sc_hd__nand4_2 _11125_ (.A(\a_h[4] ),
    .B(\a_h[5] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02068_));
 sky130_fd_sc_hd__a22o_2 _11126_ (.A1(\a_h[3] ),
    .A2(\b_h[5] ),
    .B1(_02066_),
    .B2(_02068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02069_));
 sky130_fd_sc_hd__a41o_2 _11127_ (.A1(\a_h[4] ),
    .A2(\a_h[5] ),
    .A3(\b_h[3] ),
    .A4(\b_h[4] ),
    .B1(_02063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02070_));
 sky130_fd_sc_hd__o221ai_2 _11128_ (.A1(_09406_),
    .A2(_09602_),
    .B1(_02020_),
    .B2(_02067_),
    .C1(_02066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02071_));
 sky130_fd_sc_hd__a21o_2 _11129_ (.A1(_02066_),
    .A2(_02068_),
    .B1(_02063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02072_));
 sky130_fd_sc_hd__nand2_2 _11130_ (.A(_02071_),
    .B(_02072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02073_));
 sky130_fd_sc_hd__o21ai_2 _11131_ (.A1(_02065_),
    .A2(_02070_),
    .B1(_02069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02074_));
 sky130_fd_sc_hd__o21ai_2 _11132_ (.A1(_01857_),
    .A2(_02007_),
    .B1(_02003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02075_));
 sky130_fd_sc_hd__a22o_2 _11133_ (.A1(_01962_),
    .A2(_02004_),
    .B1(_02008_),
    .B2(_02003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02076_));
 sky130_fd_sc_hd__a22oi_2 _11134_ (.A1(_01962_),
    .A2(_02004_),
    .B1(_02008_),
    .B2(_02003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_2 _11135_ (.A(\a_h[6] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_2 _11136_ (.A(\a_h[8] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02079_));
 sky130_fd_sc_hd__a22oi_2 _11137_ (.A1(\a_h[8] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_2 _11138_ (.A(_02006_),
    .B(_02079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_2 _11139_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02082_));
 sky130_fd_sc_hd__nand4_2 _11140_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02083_));
 sky130_fd_sc_hd__o2bb2ai_2 _11141_ (.A1_N(_02081_),
    .A2_N(_02083_),
    .B1(_09439_),
    .B2(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02084_));
 sky130_fd_sc_hd__nand3_2 _11142_ (.A(_02083_),
    .B(\b_h[2] ),
    .C(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02085_));
 sky130_fd_sc_hd__a21oi_2 _11143_ (.A1(_02081_),
    .A2(_02083_),
    .B1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02086_));
 sky130_fd_sc_hd__a21o_2 _11144_ (.A1(_02081_),
    .A2(_02083_),
    .B1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02087_));
 sky130_fd_sc_hd__o21a_2 _11145_ (.A1(_01857_),
    .A2(_02082_),
    .B1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02088_));
 sky130_fd_sc_hd__o21ai_2 _11146_ (.A1(_01857_),
    .A2(_02082_),
    .B1(_02078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02089_));
 sky130_fd_sc_hd__o2bb2ai_2 _11147_ (.A1_N(_02005_),
    .A2_N(_02075_),
    .B1(_02080_),
    .B2(_02089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02090_));
 sky130_fd_sc_hd__o211ai_2 _11148_ (.A1(_02080_),
    .A2(_02089_),
    .B1(_02076_),
    .C1(_02087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02091_));
 sky130_fd_sc_hd__o211ai_2 _11149_ (.A1(_02085_),
    .A2(_02080_),
    .B1(_02077_),
    .C1(_02084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02092_));
 sky130_fd_sc_hd__o21ai_2 _11150_ (.A1(_02086_),
    .A2(_02090_),
    .B1(_02092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02093_));
 sky130_fd_sc_hd__nand2_2 _11151_ (.A(_02093_),
    .B(_02073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02094_));
 sky130_fd_sc_hd__and3_2 _11152_ (.A(_02074_),
    .B(_02091_),
    .C(_02092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02095_));
 sky130_fd_sc_hd__o2111ai_2 _11153_ (.A1(_02086_),
    .A2(_02090_),
    .B1(_02092_),
    .C1(_02072_),
    .D1(_02071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02096_));
 sky130_fd_sc_hd__o211ai_2 _11154_ (.A1(_02086_),
    .A2(_02090_),
    .B1(_02092_),
    .C1(_02073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02097_));
 sky130_fd_sc_hd__a21o_2 _11155_ (.A1(_02091_),
    .A2(_02092_),
    .B1(_02073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02098_));
 sky130_fd_sc_hd__nand3_2 _11156_ (.A(_02098_),
    .B(_02061_),
    .C(_02097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_2 _11157_ (.A(_02062_),
    .B(_02094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02100_));
 sky130_fd_sc_hd__nand3_2 _11158_ (.A(_02062_),
    .B(_02094_),
    .C(_02096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02101_));
 sky130_fd_sc_hd__nand2_2 _11159_ (.A(_02099_),
    .B(_02101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02102_));
 sky130_fd_sc_hd__a21oi_2 _11160_ (.A1(_02019_),
    .A2(_02023_),
    .B1(_02021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_2 _11161_ (.A(\a_h[2] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02104_));
 sky130_fd_sc_hd__a22oi_2 _11162_ (.A1(\a_h[2] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02105_));
 sky130_fd_sc_hd__nand2_2 _11163_ (.A(_02037_),
    .B(_02104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_2 _11164_ (.A(\a_h[2] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02107_));
 sky130_fd_sc_hd__nand4_2 _11165_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_2 _11166_ (.A(\a_h[0] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02109_));
 sky130_fd_sc_hd__a22o_2 _11167_ (.A1(\a_h[0] ),
    .A2(\b_h[8] ),
    .B1(_02106_),
    .B2(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02110_));
 sky130_fd_sc_hd__a41o_2 _11168_ (.A1(\a_h[1] ),
    .A2(\a_h[2] ),
    .A3(\b_h[6] ),
    .A4(\b_h[7] ),
    .B1(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02111_));
 sky130_fd_sc_hd__o211ai_2 _11169_ (.A1(_09177_),
    .A2(_09613_),
    .B1(_02106_),
    .C1(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02112_));
 sky130_fd_sc_hd__a21o_2 _11170_ (.A1(_02106_),
    .A2(_02108_),
    .B1(_02109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02113_));
 sky130_fd_sc_hd__nand3b_2 _11171_ (.A_N(_02103_),
    .B(_02112_),
    .C(_02113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02114_));
 sky130_fd_sc_hd__o211ai_2 _11172_ (.A1(_02111_),
    .A2(_02105_),
    .B1(_02103_),
    .C1(_02110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02115_));
 sky130_fd_sc_hd__a21o_2 _11173_ (.A1(_02114_),
    .A2(_02115_),
    .B1(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02116_));
 sky130_fd_sc_hd__nand2_2 _11174_ (.A(_02114_),
    .B(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02117_));
 sky130_fd_sc_hd__nand3_2 _11175_ (.A(_02114_),
    .B(_02115_),
    .C(_02038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_2 _11176_ (.A(_02116_),
    .B(_02118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02119_));
 sky130_fd_sc_hd__a21o_2 _11177_ (.A1(_02099_),
    .A2(_02101_),
    .B1(_02119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02120_));
 sky130_fd_sc_hd__o211ai_2 _11178_ (.A1(_02095_),
    .A2(_02100_),
    .B1(_02119_),
    .C1(_02099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_2 _11179_ (.A(_02102_),
    .B(_02119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02122_));
 sky130_fd_sc_hd__nand4_2 _11180_ (.A(_02099_),
    .B(_02101_),
    .C(_02116_),
    .D(_02118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02123_));
 sky130_fd_sc_hd__a21o_2 _11181_ (.A1(_02035_),
    .A2(_02045_),
    .B1(_02033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02124_));
 sky130_fd_sc_hd__a21oi_2 _11182_ (.A1(_02035_),
    .A2(_02045_),
    .B1(_02033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02125_));
 sky130_fd_sc_hd__nand3_2 _11183_ (.A(_02120_),
    .B(_02121_),
    .C(_02125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02126_));
 sky130_fd_sc_hd__a21oi_2 _11184_ (.A1(_02120_),
    .A2(_02121_),
    .B1(_02125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02127_));
 sky130_fd_sc_hd__nand3_2 _11185_ (.A(_02122_),
    .B(_02124_),
    .C(_02123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02128_));
 sky130_fd_sc_hd__a21o_2 _11186_ (.A1(_02126_),
    .A2(_02128_),
    .B1(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02129_));
 sky130_fd_sc_hd__o211ai_2 _11187_ (.A1(_02040_),
    .A2(_02041_),
    .B1(_02126_),
    .C1(_02128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02130_));
 sky130_fd_sc_hd__o2bb2ai_2 _11188_ (.A1_N(_02126_),
    .A2_N(_02128_),
    .B1(_02040_),
    .B2(_02041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02131_));
 sky130_fd_sc_hd__a31oi_2 _11189_ (.A1(_02120_),
    .A2(_02121_),
    .A3(_02125_),
    .B1(_02043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02132_));
 sky130_fd_sc_hd__nand3_2 _11190_ (.A(_02126_),
    .B(_02128_),
    .C(_02042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02133_));
 sky130_fd_sc_hd__o2bb2ai_2 _11191_ (.A1_N(_01984_),
    .A2_N(_02053_),
    .B1(_02051_),
    .B2(_02049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02134_));
 sky130_fd_sc_hd__a21boi_2 _11192_ (.A1(_02053_),
    .A2(_01984_),
    .B1_N(_02052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02135_));
 sky130_fd_sc_hd__and3_2 _11193_ (.A(_02129_),
    .B(_02130_),
    .C(_02135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02136_));
 sky130_fd_sc_hd__nand3_2 _11194_ (.A(_02129_),
    .B(_02130_),
    .C(_02135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02137_));
 sky130_fd_sc_hd__o31ai_2 _11195_ (.A1(_01991_),
    .A2(_02055_),
    .A3(_02056_),
    .B1(_01990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_2 _11196_ (.A(_02136_),
    .B(_02138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02139_));
 sky130_fd_sc_hd__a22oi_2 _11197_ (.A1(_02132_),
    .A2(_02128_),
    .B1(_02054_),
    .B2(_02052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02140_));
 sky130_fd_sc_hd__nand3_2 _11198_ (.A(_02131_),
    .B(_02134_),
    .C(_02133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_2 _11199_ (.A(_02137_),
    .B(_02141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02142_));
 sky130_fd_sc_hd__o211a_2 _11200_ (.A1(_02055_),
    .A2(_02056_),
    .B1(_01991_),
    .C1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02143_));
 sky130_fd_sc_hd__o211ai_2 _11201_ (.A1(_02055_),
    .A2(_02056_),
    .B1(_01991_),
    .C1(_02137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02144_));
 sky130_fd_sc_hd__a311o_2 _11202_ (.A1(_02060_),
    .A2(_02138_),
    .A3(_02142_),
    .B1(_02143_),
    .C1(_02139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02145_));
 sky130_fd_sc_hd__o211ai_2 _11203_ (.A1(_02055_),
    .A2(_02056_),
    .B1(_01992_),
    .C1(_01993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02146_));
 sky130_fd_sc_hd__a31oi_2 _11204_ (.A1(_02060_),
    .A2(_02138_),
    .A3(_02142_),
    .B1(_02146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02147_));
 sky130_fd_sc_hd__a211oi_2 _11205_ (.A1(_02145_),
    .A2(_02146_),
    .B1(_02147_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00282_));
 sky130_fd_sc_hd__nor2_2 _11206_ (.A(_02139_),
    .B(_02147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02148_));
 sky130_fd_sc_hd__a21oi_2 _11207_ (.A1(_02042_),
    .A2(_02126_),
    .B1(_02127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02149_));
 sky130_fd_sc_hd__o2bb2ai_2 _11208_ (.A1_N(_02099_),
    .A2_N(_02119_),
    .B1(_02100_),
    .B2(_02095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02150_));
 sky130_fd_sc_hd__a21boi_2 _11209_ (.A1(_02099_),
    .A2(_02119_),
    .B1_N(_02101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02151_));
 sky130_fd_sc_hd__a2bb2oi_2 _11210_ (.A1_N(_02086_),
    .A2_N(_02090_),
    .B1(_02092_),
    .B2(_02074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02152_));
 sky130_fd_sc_hd__a21boi_2 _11211_ (.A1(_02073_),
    .A2(_02091_),
    .B1_N(_02092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02153_));
 sky130_fd_sc_hd__and2_2 _11212_ (.A(\a_h[4] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02154_));
 sky130_fd_sc_hd__nand2_2 _11213_ (.A(\a_h[4] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_2 _11214_ (.A(\a_h[6] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02156_));
 sky130_fd_sc_hd__a22oi_2 _11215_ (.A1(\a_h[6] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_2 _11216_ (.A(_02067_),
    .B(_02156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_2 _11217_ (.A(\a_h[6] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02159_));
 sky130_fd_sc_hd__nand4_2 _11218_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02160_));
 sky130_fd_sc_hd__a21oi_2 _11219_ (.A1(_02158_),
    .A2(_02160_),
    .B1(_02154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02161_));
 sky130_fd_sc_hd__o211a_2 _11220_ (.A1(_02064_),
    .A2(_02159_),
    .B1(_02154_),
    .C1(_02158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02162_));
 sky130_fd_sc_hd__nor2_2 _11221_ (.A(_02161_),
    .B(_02162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02163_));
 sky130_fd_sc_hd__o21ai_2 _11222_ (.A1(_02078_),
    .A2(_02080_),
    .B1(_02083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02164_));
 sky130_fd_sc_hd__nand2_2 _11223_ (.A(\a_h[7] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2_2 _11224_ (.A(\a_h[8] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02166_));
 sky130_fd_sc_hd__nand2_2 _11225_ (.A(\a_h[9] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02167_));
 sky130_fd_sc_hd__a22oi_2 _11226_ (.A1(\a_h[9] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_2 _11227_ (.A(_02166_),
    .B(_02167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02169_));
 sky130_fd_sc_hd__nand2_2 _11228_ (.A(\a_h[9] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02170_));
 sky130_fd_sc_hd__nand4_2 _11229_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02171_));
 sky130_fd_sc_hd__o221ai_2 _11230_ (.A1(_09449_),
    .A2(_09592_),
    .B1(_02079_),
    .B2(_02170_),
    .C1(_02169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02172_));
 sky130_fd_sc_hd__a21o_2 _11231_ (.A1(_02169_),
    .A2(_02171_),
    .B1(_02165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02173_));
 sky130_fd_sc_hd__o2111ai_2 _11232_ (.A1(_02079_),
    .A2(_02170_),
    .B1(\a_h[7] ),
    .C1(\b_h[2] ),
    .D1(_02169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02174_));
 sky130_fd_sc_hd__a22o_2 _11233_ (.A1(\a_h[7] ),
    .A2(\b_h[2] ),
    .B1(_02169_),
    .B2(_02171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02175_));
 sky130_fd_sc_hd__nand3_2 _11234_ (.A(_02175_),
    .B(_02164_),
    .C(_02174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02176_));
 sky130_fd_sc_hd__o211ai_2 _11235_ (.A1(_02080_),
    .A2(_02088_),
    .B1(_02172_),
    .C1(_02173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_2 _11236_ (.A(_02176_),
    .B(_02177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_2 _11237_ (.A(_02177_),
    .B(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02179_));
 sky130_fd_sc_hd__nand3_2 _11238_ (.A(_02176_),
    .B(_02177_),
    .C(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02180_));
 sky130_fd_sc_hd__o21ai_2 _11239_ (.A1(_02161_),
    .A2(_02162_),
    .B1(_02178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_2 _11240_ (.A(_02178_),
    .B(_02163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02182_));
 sky130_fd_sc_hd__o211ai_2 _11241_ (.A1(_02161_),
    .A2(_02162_),
    .B1(_02176_),
    .C1(_02177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02183_));
 sky130_fd_sc_hd__a21oi_2 _11242_ (.A1(_02182_),
    .A2(_02183_),
    .B1(_02153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02184_));
 sky130_fd_sc_hd__nand3_2 _11243_ (.A(_02181_),
    .B(_02152_),
    .C(_02180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02185_));
 sky130_fd_sc_hd__nand3_2 _11244_ (.A(_02153_),
    .B(_02182_),
    .C(_02183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02186_));
 sky130_fd_sc_hd__a21o_2 _11245_ (.A1(_02063_),
    .A2(_02068_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02187_));
 sky130_fd_sc_hd__a21oi_2 _11246_ (.A1(_02063_),
    .A2(_02068_),
    .B1(_02065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_2 _11247_ (.A(\a_h[1] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02189_));
 sky130_fd_sc_hd__nand2_2 _11248_ (.A(\a_h[3] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02190_));
 sky130_fd_sc_hd__a22oi_2 _11249_ (.A1(\a_h[3] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02191_));
 sky130_fd_sc_hd__nand2_2 _11250_ (.A(_02107_),
    .B(_02190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_2 _11251_ (.A(\a_h[3] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02193_));
 sky130_fd_sc_hd__nand4_2 _11252_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02194_));
 sky130_fd_sc_hd__a22o_2 _11253_ (.A1(\a_h[1] ),
    .A2(\b_h[8] ),
    .B1(_02192_),
    .B2(_02194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02195_));
 sky130_fd_sc_hd__a41o_2 _11254_ (.A1(\a_h[2] ),
    .A2(\a_h[3] ),
    .A3(\b_h[6] ),
    .A4(\b_h[7] ),
    .B1(_02189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02196_));
 sky130_fd_sc_hd__o21ai_2 _11255_ (.A1(_02104_),
    .A2(_02193_),
    .B1(_02189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02197_));
 sky130_fd_sc_hd__a21o_2 _11256_ (.A1(_02192_),
    .A2(_02194_),
    .B1(_02189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02198_));
 sky130_fd_sc_hd__o211ai_2 _11257_ (.A1(_02191_),
    .A2(_02197_),
    .B1(_02187_),
    .C1(_02198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02199_));
 sky130_fd_sc_hd__o211ai_2 _11258_ (.A1(_02196_),
    .A2(_02191_),
    .B1(_02188_),
    .C1(_02195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02200_));
 sky130_fd_sc_hd__o21a_2 _11259_ (.A1(_09177_),
    .A2(_09613_),
    .B1(_02108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02201_));
 sky130_fd_sc_hd__a21oi_2 _11260_ (.A1(_02108_),
    .A2(_02109_),
    .B1(_02105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02202_));
 sky130_fd_sc_hd__o2bb2a_2 _11261_ (.A1_N(_02199_),
    .A2_N(_02200_),
    .B1(_02201_),
    .B2(_02105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02203_));
 sky130_fd_sc_hd__o2bb2ai_2 _11262_ (.A1_N(_02199_),
    .A2_N(_02200_),
    .B1(_02201_),
    .B2(_02105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_2 _11263_ (.A(_02199_),
    .B(_02202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02205_));
 sky130_fd_sc_hd__and3_2 _11264_ (.A(_02199_),
    .B(_02200_),
    .C(_02202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02206_));
 sky130_fd_sc_hd__nand3_2 _11265_ (.A(_02199_),
    .B(_02200_),
    .C(_02202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02207_));
 sky130_fd_sc_hd__a221oi_2 _11266_ (.A1(_02108_),
    .A2(_02109_),
    .B1(_02199_),
    .B2(_02200_),
    .C1(_02105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02208_));
 sky130_fd_sc_hd__a21bo_2 _11267_ (.A1(_02199_),
    .A2(_02200_),
    .B1_N(_02202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02209_));
 sky130_fd_sc_hd__o211a_2 _11268_ (.A1(_02105_),
    .A2(_02201_),
    .B1(_02200_),
    .C1(_02199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02210_));
 sky130_fd_sc_hd__o211ai_2 _11269_ (.A1(_02105_),
    .A2(_02201_),
    .B1(_02200_),
    .C1(_02199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02211_));
 sky130_fd_sc_hd__nand2_2 _11270_ (.A(_02209_),
    .B(_02211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2_2 _11271_ (.A(_02204_),
    .B(_02207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02213_));
 sky130_fd_sc_hd__nand4_2 _11272_ (.A(_02185_),
    .B(_02186_),
    .C(_02209_),
    .D(_02211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02214_));
 sky130_fd_sc_hd__o2bb2ai_2 _11273_ (.A1_N(_02185_),
    .A2_N(_02186_),
    .B1(_02208_),
    .B2(_02210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02215_));
 sky130_fd_sc_hd__nand3_2 _11274_ (.A(_02215_),
    .B(_02150_),
    .C(_02214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02216_));
 sky130_fd_sc_hd__nand4_2 _11275_ (.A(_02185_),
    .B(_02186_),
    .C(_02204_),
    .D(_02207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02217_));
 sky130_fd_sc_hd__o2bb2ai_2 _11276_ (.A1_N(_02185_),
    .A2_N(_02186_),
    .B1(_02203_),
    .B2(_02206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02218_));
 sky130_fd_sc_hd__nand3_2 _11277_ (.A(_02151_),
    .B(_02217_),
    .C(_02218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2_2 _11278_ (.A(\a_h[0] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02220_));
 sky130_fd_sc_hd__and2_2 _11279_ (.A(_02115_),
    .B(_02117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02221_));
 sky130_fd_sc_hd__and3_2 _11280_ (.A(_02115_),
    .B(_02117_),
    .C(_02220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02222_));
 sky130_fd_sc_hd__a21oi_2 _11281_ (.A1(_02115_),
    .A2(_02117_),
    .B1(_02220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_2 _11282_ (.A(_02222_),
    .B(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02224_));
 sky130_fd_sc_hd__inv_2 _11283_ (.A(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02225_));
 sky130_fd_sc_hd__nand3_2 _11284_ (.A(_02216_),
    .B(_02219_),
    .C(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02226_));
 sky130_fd_sc_hd__o2bb2ai_2 _11285_ (.A1_N(_02216_),
    .A2_N(_02219_),
    .B1(_02222_),
    .B2(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02227_));
 sky130_fd_sc_hd__o211ai_2 _11286_ (.A1(_02222_),
    .A2(_02223_),
    .B1(_02216_),
    .C1(_02219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02228_));
 sky130_fd_sc_hd__a21o_2 _11287_ (.A1(_02216_),
    .A2(_02219_),
    .B1(_02225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02229_));
 sky130_fd_sc_hd__o211a_2 _11288_ (.A1(_02127_),
    .A2(_02132_),
    .B1(_02226_),
    .C1(_02227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02230_));
 sky130_fd_sc_hd__o211ai_2 _11289_ (.A1(_02127_),
    .A2(_02132_),
    .B1(_02226_),
    .C1(_02227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02231_));
 sky130_fd_sc_hd__nand3_2 _11290_ (.A(_02229_),
    .B(_02149_),
    .C(_02228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02232_));
 sky130_fd_sc_hd__nand2_2 _11291_ (.A(_02231_),
    .B(_02232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02233_));
 sky130_fd_sc_hd__a22oi_2 _11292_ (.A1(_02140_),
    .A2(_02131_),
    .B1(_02232_),
    .B2(_02231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02234_));
 sky130_fd_sc_hd__a31oi_2 _11293_ (.A1(_02149_),
    .A2(_02228_),
    .A3(_02229_),
    .B1(_02141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02235_));
 sky130_fd_sc_hd__a21oi_2 _11294_ (.A1(_02235_),
    .A2(_02231_),
    .B1(_02234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02236_));
 sky130_fd_sc_hd__xor2_2 _11295_ (.A(_02144_),
    .B(_02236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02237_));
 sky130_fd_sc_hd__a21oi_2 _11296_ (.A1(_02237_),
    .A2(_02148_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02238_));
 sky130_fd_sc_hd__o21a_2 _11297_ (.A1(_02148_),
    .A2(_02237_),
    .B1(_02238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00283_));
 sky130_fd_sc_hd__a31o_2 _11298_ (.A1(_02151_),
    .A2(_02217_),
    .A3(_02218_),
    .B1(_02224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02239_));
 sky130_fd_sc_hd__nand2_2 _11299_ (.A(_02216_),
    .B(_02239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02240_));
 sky130_fd_sc_hd__a21boi_2 _11300_ (.A1(_02219_),
    .A2(_02225_),
    .B1_N(_02216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02241_));
 sky130_fd_sc_hd__o2bb2a_2 _11301_ (.A1_N(\a_h[1] ),
    .A2_N(\b_h[9] ),
    .B1(_09635_),
    .B2(_09177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02242_));
 sky130_fd_sc_hd__and4_2 _11302_ (.A(\a_h[0] ),
    .B(\a_h[1] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02243_));
 sky130_fd_sc_hd__or2_2 _11303_ (.A(_02242_),
    .B(_02243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02244_));
 sky130_fd_sc_hd__and2_2 _11304_ (.A(_02200_),
    .B(_02205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02245_));
 sky130_fd_sc_hd__o21ai_2 _11305_ (.A1(_02242_),
    .A2(_02243_),
    .B1(_02245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02246_));
 sky130_fd_sc_hd__a211o_2 _11306_ (.A1(_02200_),
    .A2(_02205_),
    .B1(_02242_),
    .C1(_02243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02247_));
 sky130_fd_sc_hd__and2_2 _11307_ (.A(_02246_),
    .B(_02247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02248_));
 sky130_fd_sc_hd__nand2_2 _11308_ (.A(_02246_),
    .B(_02247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02249_));
 sky130_fd_sc_hd__a31oi_2 _11309_ (.A1(_02153_),
    .A2(_02182_),
    .A3(_02183_),
    .B1(_02213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02250_));
 sky130_fd_sc_hd__a21oi_2 _11310_ (.A1(_02186_),
    .A2(_02212_),
    .B1(_02184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02251_));
 sky130_fd_sc_hd__a21o_2 _11311_ (.A1(_02155_),
    .A2(_02160_),
    .B1(_02157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02252_));
 sky130_fd_sc_hd__a21oi_2 _11312_ (.A1(_02155_),
    .A2(_02160_),
    .B1(_02157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_2 _11313_ (.A(\a_h[2] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02254_));
 sky130_fd_sc_hd__nand2_2 _11314_ (.A(\a_h[4] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_2 _11315_ (.A(\a_h[4] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02256_));
 sky130_fd_sc_hd__nand4_2 _11316_ (.A(\a_h[3] ),
    .B(\a_h[4] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02257_));
 sky130_fd_sc_hd__nand2_2 _11317_ (.A(_02193_),
    .B(_02256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02258_));
 sky130_fd_sc_hd__o2bb2ai_2 _11318_ (.A1_N(_02257_),
    .A2_N(_02258_),
    .B1(_09395_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02259_));
 sky130_fd_sc_hd__o2111ai_2 _11319_ (.A1(_02190_),
    .A2(_02255_),
    .B1(\a_h[2] ),
    .C1(\b_h[8] ),
    .D1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02260_));
 sky130_fd_sc_hd__a21o_2 _11320_ (.A1(_02257_),
    .A2(_02258_),
    .B1(_02254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02261_));
 sky130_fd_sc_hd__o221ai_2 _11321_ (.A1(_09395_),
    .A2(_09613_),
    .B1(_02190_),
    .B2(_02255_),
    .C1(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02262_));
 sky130_fd_sc_hd__nand3_2 _11322_ (.A(_02253_),
    .B(_02259_),
    .C(_02260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02263_));
 sky130_fd_sc_hd__nand3_2 _11323_ (.A(_02261_),
    .B(_02262_),
    .C(_02252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02264_));
 sky130_fd_sc_hd__a21oi_2 _11324_ (.A1(_02189_),
    .A2(_02194_),
    .B1(_02191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02265_));
 sky130_fd_sc_hd__nand3b_2 _11325_ (.A_N(_02265_),
    .B(_02264_),
    .C(_02263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02266_));
 sky130_fd_sc_hd__a21bo_2 _11326_ (.A1(_02263_),
    .A2(_02264_),
    .B1_N(_02265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02267_));
 sky130_fd_sc_hd__a22o_2 _11327_ (.A1(_02192_),
    .A2(_02197_),
    .B1(_02263_),
    .B2(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02268_));
 sky130_fd_sc_hd__nand4_2 _11328_ (.A(_02192_),
    .B(_02197_),
    .C(_02263_),
    .D(_02264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_2 _11329_ (.A(_02268_),
    .B(_02269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_2 _11330_ (.A(_02266_),
    .B(_02267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02271_));
 sky130_fd_sc_hd__nand2_2 _11331_ (.A(_02176_),
    .B(_02179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02272_));
 sky130_fd_sc_hd__a21boi_2 _11332_ (.A1(_02163_),
    .A2(_02177_),
    .B1_N(_02176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02273_));
 sky130_fd_sc_hd__nand2_2 _11333_ (.A(\a_h[8] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_2 _11334_ (.A(\a_h[10] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02275_));
 sky130_fd_sc_hd__a22oi_2 _11335_ (.A1(\a_h[10] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02276_));
 sky130_fd_sc_hd__nand2_2 _11336_ (.A(_02170_),
    .B(_02275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_2 _11337_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02278_));
 sky130_fd_sc_hd__nand4_2 _11338_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02279_));
 sky130_fd_sc_hd__o2bb2ai_2 _11339_ (.A1_N(_02277_),
    .A2_N(_02279_),
    .B1(_09460_),
    .B2(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02280_));
 sky130_fd_sc_hd__o2111ai_2 _11340_ (.A1(_01857_),
    .A2(_02278_),
    .B1(\a_h[8] ),
    .C1(\b_h[2] ),
    .D1(_02277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02281_));
 sky130_fd_sc_hd__a21o_2 _11341_ (.A1(_02277_),
    .A2(_02279_),
    .B1(_02274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02282_));
 sky130_fd_sc_hd__o22a_2 _11342_ (.A1(_09460_),
    .A2(_09592_),
    .B1(_01857_),
    .B2(_02278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02283_));
 sky130_fd_sc_hd__o221ai_2 _11343_ (.A1(_09460_),
    .A2(_09592_),
    .B1(_01857_),
    .B2(_02278_),
    .C1(_02277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02284_));
 sky130_fd_sc_hd__nand2_2 _11344_ (.A(_02165_),
    .B(_02171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02285_));
 sky130_fd_sc_hd__o21ai_2 _11345_ (.A1(_02165_),
    .A2(_02168_),
    .B1(_02171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_2 _11346_ (.A(_02169_),
    .B(_02285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02287_));
 sky130_fd_sc_hd__nand3_2 _11347_ (.A(_02282_),
    .B(_02284_),
    .C(_02287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02288_));
 sky130_fd_sc_hd__nand3_2 _11348_ (.A(_02280_),
    .B(_02281_),
    .C(_02286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_2 _11349_ (.A(_02288_),
    .B(_02289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_2 _11350_ (.A(\a_h[5] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02291_));
 sky130_fd_sc_hd__nand2_2 _11351_ (.A(\a_h[7] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_2 _11352_ (.A(\a_h[7] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02293_));
 sky130_fd_sc_hd__and4_2 _11353_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02294_));
 sky130_fd_sc_hd__nand4_2 _11354_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_2 _11355_ (.A(_02159_),
    .B(_02293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02296_));
 sky130_fd_sc_hd__a22oi_2 _11356_ (.A1(\a_h[5] ),
    .A2(\b_h[5] ),
    .B1(_02295_),
    .B2(_02296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02297_));
 sky130_fd_sc_hd__o2bb2ai_2 _11357_ (.A1_N(_02295_),
    .A2_N(_02296_),
    .B1(_09428_),
    .B2(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02298_));
 sky130_fd_sc_hd__a21oi_2 _11358_ (.A1(_02159_),
    .A2(_02293_),
    .B1(_02291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02299_));
 sky130_fd_sc_hd__o21ai_2 _11359_ (.A1(_02156_),
    .A2(_02292_),
    .B1(_02299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02300_));
 sky130_fd_sc_hd__a21oi_2 _11360_ (.A1(_02295_),
    .A2(_02299_),
    .B1(_02297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02301_));
 sky130_fd_sc_hd__nand2_2 _11361_ (.A(_02298_),
    .B(_02300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02302_));
 sky130_fd_sc_hd__nand2_2 _11362_ (.A(_02290_),
    .B(_02301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02303_));
 sky130_fd_sc_hd__nand3_2 _11363_ (.A(_02288_),
    .B(_02289_),
    .C(_02302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02304_));
 sky130_fd_sc_hd__a21oi_2 _11364_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02305_));
 sky130_fd_sc_hd__a21o_2 _11365_ (.A1(_02288_),
    .A2(_02289_),
    .B1(_02301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02306_));
 sky130_fd_sc_hd__nand4_2 _11366_ (.A(_02288_),
    .B(_02289_),
    .C(_02298_),
    .D(_02300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02307_));
 sky130_fd_sc_hd__a21oi_2 _11367_ (.A1(_02176_),
    .A2(_02179_),
    .B1(_02305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02308_));
 sky130_fd_sc_hd__nand3_2 _11368_ (.A(_02272_),
    .B(_02306_),
    .C(_02307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02309_));
 sky130_fd_sc_hd__nand3_2 _11369_ (.A(_02273_),
    .B(_02303_),
    .C(_02304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02310_));
 sky130_fd_sc_hd__nand4_2 _11370_ (.A(_02266_),
    .B(_02267_),
    .C(_02309_),
    .D(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02311_));
 sky130_fd_sc_hd__a22o_2 _11371_ (.A1(_02266_),
    .A2(_02267_),
    .B1(_02309_),
    .B2(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02312_));
 sky130_fd_sc_hd__nand4_2 _11372_ (.A(_02268_),
    .B(_02269_),
    .C(_02309_),
    .D(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02313_));
 sky130_fd_sc_hd__a22o_2 _11373_ (.A1(_02268_),
    .A2(_02269_),
    .B1(_02309_),
    .B2(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02314_));
 sky130_fd_sc_hd__o211ai_2 _11374_ (.A1(_02184_),
    .A2(_02250_),
    .B1(_02313_),
    .C1(_02314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02315_));
 sky130_fd_sc_hd__nand3_2 _11375_ (.A(_02312_),
    .B(_02251_),
    .C(_02311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02316_));
 sky130_fd_sc_hd__nand4_2 _11376_ (.A(_02246_),
    .B(_02247_),
    .C(_02315_),
    .D(_02316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02317_));
 sky130_fd_sc_hd__a22o_2 _11377_ (.A1(_02246_),
    .A2(_02247_),
    .B1(_02315_),
    .B2(_02316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02318_));
 sky130_fd_sc_hd__a21o_2 _11378_ (.A1(_02315_),
    .A2(_02316_),
    .B1(_02249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02319_));
 sky130_fd_sc_hd__nand3_2 _11379_ (.A(_02249_),
    .B(_02315_),
    .C(_02316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02320_));
 sky130_fd_sc_hd__a21oi_2 _11380_ (.A1(_02319_),
    .A2(_02320_),
    .B1(_02240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02321_));
 sky130_fd_sc_hd__nand3_2 _11381_ (.A(_02241_),
    .B(_02317_),
    .C(_02318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02322_));
 sky130_fd_sc_hd__nand3_2 _11382_ (.A(_02240_),
    .B(_02319_),
    .C(_02320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02323_));
 sky130_fd_sc_hd__o2bb2ai_2 _11383_ (.A1_N(_02322_),
    .A2_N(_02323_),
    .B1(_02220_),
    .B2(_02221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_2 _11384_ (.A(_02323_),
    .B(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02325_));
 sky130_fd_sc_hd__a21bo_2 _11385_ (.A1(_02322_),
    .A2(_02323_),
    .B1_N(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02326_));
 sky130_fd_sc_hd__a31o_2 _11386_ (.A1(_02240_),
    .A2(_02319_),
    .A3(_02320_),
    .B1(_02223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02327_));
 sky130_fd_sc_hd__o21ai_2 _11387_ (.A1(_02321_),
    .A2(_02325_),
    .B1(_02324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02328_));
 sky130_fd_sc_hd__a31oi_2 _11388_ (.A1(_02131_),
    .A2(_02232_),
    .A3(_02140_),
    .B1(_02230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02329_));
 sky130_fd_sc_hd__o211ai_2 _11389_ (.A1(_02321_),
    .A2(_02327_),
    .B1(_02329_),
    .C1(_02326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02330_));
 sky130_fd_sc_hd__o221ai_2 _11390_ (.A1(_02321_),
    .A2(_02325_),
    .B1(_02230_),
    .B2(_02235_),
    .C1(_02324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02331_));
 sky130_fd_sc_hd__nand2_2 _11391_ (.A(_02330_),
    .B(_02331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02332_));
 sky130_fd_sc_hd__o22ai_2 _11392_ (.A1(_02136_),
    .A2(_02138_),
    .B1(_02144_),
    .B2(_02234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02333_));
 sky130_fd_sc_hd__o22ai_2 _11393_ (.A1(_02143_),
    .A2(_02236_),
    .B1(_02333_),
    .B2(_02147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02334_));
 sky130_fd_sc_hd__a21o_2 _11394_ (.A1(_02334_),
    .A2(_02332_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02335_));
 sky130_fd_sc_hd__o21ba_2 _11395_ (.A1(_02332_),
    .A2(_02334_),
    .B1_N(_02335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00284_));
 sky130_fd_sc_hd__a32oi_2 _11396_ (.A1(_02251_),
    .A2(_02311_),
    .A3(_02312_),
    .B1(_02315_),
    .B2(_02249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02336_));
 sky130_fd_sc_hd__a21boi_2 _11397_ (.A1(_02248_),
    .A2(_02316_),
    .B1_N(_02315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02337_));
 sky130_fd_sc_hd__nand2_2 _11398_ (.A(\b_h[9] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02338_));
 sky130_fd_sc_hd__and4_2 _11399_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02339_));
 sky130_fd_sc_hd__nand4_2 _11400_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02340_));
 sky130_fd_sc_hd__a22oi_2 _11401_ (.A1(\a_h[2] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02341_));
 sky130_fd_sc_hd__nand2_2 _11402_ (.A(\a_h[0] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02342_));
 sky130_fd_sc_hd__o22a_2 _11403_ (.A1(_09177_),
    .A2(_09646_),
    .B1(_02339_),
    .B2(_02341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02343_));
 sky130_fd_sc_hd__and4b_2 _11404_ (.A_N(_02341_),
    .B(\b_h[11] ),
    .C(\a_h[0] ),
    .D(_02340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02344_));
 sky130_fd_sc_hd__nor2_2 _11405_ (.A(_02343_),
    .B(_02344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02345_));
 sky130_fd_sc_hd__o32ai_2 _11406_ (.A1(_09624_),
    .A2(_09635_),
    .A3(_01855_),
    .B1(_02343_),
    .B2(_02344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02346_));
 sky130_fd_sc_hd__nand2_2 _11407_ (.A(_02243_),
    .B(_02345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_2 _11408_ (.A(_02346_),
    .B(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02348_));
 sky130_fd_sc_hd__a21bo_2 _11409_ (.A1(_02264_),
    .A2(_02265_),
    .B1_N(_02263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02349_));
 sky130_fd_sc_hd__inv_2 _11410_ (.A(_02349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02350_));
 sky130_fd_sc_hd__and3_2 _11411_ (.A(_02349_),
    .B(_02347_),
    .C(_02346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02351_));
 sky130_fd_sc_hd__inv_2 _11412_ (.A(_02351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02352_));
 sky130_fd_sc_hd__a21oi_2 _11413_ (.A1(_02346_),
    .A2(_02347_),
    .B1(_02349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_2 _11414_ (.A(_02351_),
    .B(_02353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02354_));
 sky130_fd_sc_hd__o22ai_2 _11415_ (.A1(_01857_),
    .A2(_02278_),
    .B1(_02274_),
    .B2(_02276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02355_));
 sky130_fd_sc_hd__and2_2 _11416_ (.A(\a_h[9] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02356_));
 sky130_fd_sc_hd__nand2_2 _11417_ (.A(\a_h[9] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_2 _11418_ (.A(\a_h[10] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02358_));
 sky130_fd_sc_hd__nand2_2 _11419_ (.A(\a_h[11] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02359_));
 sky130_fd_sc_hd__a22oi_2 _11420_ (.A1(\a_h[11] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_2 _11421_ (.A(_02358_),
    .B(_02359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_2 _11422_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02362_));
 sky130_fd_sc_hd__nand3_2 _11423_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02363_));
 sky130_fd_sc_hd__nand4_2 _11424_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02364_));
 sky130_fd_sc_hd__a21oi_2 _11425_ (.A1(_02361_),
    .A2(_02364_),
    .B1(_02356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02365_));
 sky130_fd_sc_hd__a21o_2 _11426_ (.A1(_02361_),
    .A2(_02364_),
    .B1(_02356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02366_));
 sky130_fd_sc_hd__o211a_2 _11427_ (.A1(_09526_),
    .A2(_02363_),
    .B1(_02356_),
    .C1(_02361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02367_));
 sky130_fd_sc_hd__o2111ai_2 _11428_ (.A1(_09526_),
    .A2(_02363_),
    .B1(\b_h[2] ),
    .C1(\a_h[9] ),
    .D1(_02361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02368_));
 sky130_fd_sc_hd__a21oi_2 _11429_ (.A1(_02366_),
    .A2(_02368_),
    .B1(_02355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02369_));
 sky130_fd_sc_hd__o22ai_2 _11430_ (.A1(_02276_),
    .A2(_02283_),
    .B1(_02365_),
    .B2(_02367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_2 _11431_ (.A(_02366_),
    .B(_02355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02371_));
 sky130_fd_sc_hd__nand3_2 _11432_ (.A(_02366_),
    .B(_02368_),
    .C(_02355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_2 _11433_ (.A(\a_h[6] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_2 _11434_ (.A(\a_h[8] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02374_));
 sky130_fd_sc_hd__a22oi_2 _11435_ (.A1(\a_h[8] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_2 _11436_ (.A(_02292_),
    .B(_02374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02376_));
 sky130_fd_sc_hd__nand4_2 _11437_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02377_));
 sky130_fd_sc_hd__o2bb2a_2 _11438_ (.A1_N(_02376_),
    .A2_N(_02377_),
    .B1(_09439_),
    .B2(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02378_));
 sky130_fd_sc_hd__a22o_2 _11439_ (.A1(\a_h[6] ),
    .A2(\b_h[5] ),
    .B1(_02376_),
    .B2(_02377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02379_));
 sky130_fd_sc_hd__and4_2 _11440_ (.A(_02376_),
    .B(_02377_),
    .C(\a_h[6] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02380_));
 sky130_fd_sc_hd__nand4_2 _11441_ (.A(_02376_),
    .B(_02377_),
    .C(\a_h[6] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_2 _11442_ (.A(_02379_),
    .B(_02381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02382_));
 sky130_fd_sc_hd__a21o_2 _11443_ (.A1(_02370_),
    .A2(_02372_),
    .B1(_02382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02383_));
 sky130_fd_sc_hd__o221ai_2 _11444_ (.A1(_02378_),
    .A2(_02380_),
    .B1(_02367_),
    .B2(_02371_),
    .C1(_02370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02384_));
 sky130_fd_sc_hd__o2bb2ai_2 _11445_ (.A1_N(_02370_),
    .A2_N(_02372_),
    .B1(_02378_),
    .B2(_02380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02385_));
 sky130_fd_sc_hd__nand4_2 _11446_ (.A(_02370_),
    .B(_02372_),
    .C(_02379_),
    .D(_02381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02386_));
 sky130_fd_sc_hd__a32oi_2 _11447_ (.A1(_02282_),
    .A2(_02284_),
    .A3(_02287_),
    .B1(_02289_),
    .B2(_02302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02387_));
 sky130_fd_sc_hd__a21boi_2 _11448_ (.A1(_02301_),
    .A2(_02288_),
    .B1_N(_02289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02388_));
 sky130_fd_sc_hd__nand3_2 _11449_ (.A(_02383_),
    .B(_02384_),
    .C(_02388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02389_));
 sky130_fd_sc_hd__nand3_2 _11450_ (.A(_02385_),
    .B(_02386_),
    .C(_02387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_2 _11451_ (.A(_02291_),
    .B(_02295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_2 _11452_ (.A(_02296_),
    .B(_02391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02392_));
 sky130_fd_sc_hd__and2_2 _11453_ (.A(\a_h[3] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02393_));
 sky130_fd_sc_hd__nand2_2 _11454_ (.A(\a_h[3] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02394_));
 sky130_fd_sc_hd__nand2_2 _11455_ (.A(\a_h[5] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_2 _11456_ (.A(_02255_),
    .B(_02395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_2 _11457_ (.A(\a_h[5] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02397_));
 sky130_fd_sc_hd__and4_2 _11458_ (.A(\a_h[4] ),
    .B(\a_h[5] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02398_));
 sky130_fd_sc_hd__nand4_2 _11459_ (.A(\a_h[4] ),
    .B(\a_h[5] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02399_));
 sky130_fd_sc_hd__o221ai_2 _11460_ (.A1(_09406_),
    .A2(_09613_),
    .B1(_02256_),
    .B2(_02397_),
    .C1(_02396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02400_));
 sky130_fd_sc_hd__a21o_2 _11461_ (.A1(_02396_),
    .A2(_02399_),
    .B1(_02394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02401_));
 sky130_fd_sc_hd__o211ai_2 _11462_ (.A1(_02256_),
    .A2(_02397_),
    .B1(_02393_),
    .C1(_02396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3_2 _11463_ (.A(_02255_),
    .B(\b_h[6] ),
    .C(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02403_));
 sky130_fd_sc_hd__nand3_2 _11464_ (.A(_02395_),
    .B(\b_h[7] ),
    .C(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02404_));
 sky130_fd_sc_hd__o211ai_2 _11465_ (.A1(_09406_),
    .A2(_09613_),
    .B1(_02403_),
    .C1(_02404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_2 _11466_ (.A(_02402_),
    .B(_02405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3_2 _11467_ (.A(_02401_),
    .B(_02392_),
    .C(_02400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02407_));
 sky130_fd_sc_hd__o211ai_2 _11468_ (.A1(_02294_),
    .A2(_02299_),
    .B1(_02402_),
    .C1(_02405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02408_));
 sky130_fd_sc_hd__a21boi_2 _11469_ (.A1(_02254_),
    .A2(_02257_),
    .B1_N(_02258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02409_));
 sky130_fd_sc_hd__inv_2 _11470_ (.A(_02409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02410_));
 sky130_fd_sc_hd__a21o_2 _11471_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_2 _11472_ (.A(_02407_),
    .B(_02409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02412_));
 sky130_fd_sc_hd__nand3_2 _11473_ (.A(_02407_),
    .B(_02408_),
    .C(_02409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02413_));
 sky130_fd_sc_hd__a21oi_2 _11474_ (.A1(_02407_),
    .A2(_02408_),
    .B1(_02410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02414_));
 sky130_fd_sc_hd__and3_2 _11475_ (.A(_02407_),
    .B(_02410_),
    .C(_02408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02415_));
 sky130_fd_sc_hd__nand2_2 _11476_ (.A(_02411_),
    .B(_02413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02416_));
 sky130_fd_sc_hd__o2bb2ai_2 _11477_ (.A1_N(_02389_),
    .A2_N(_02390_),
    .B1(_02414_),
    .B2(_02415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02417_));
 sky130_fd_sc_hd__nand3_2 _11478_ (.A(_02389_),
    .B(_02390_),
    .C(_02416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02418_));
 sky130_fd_sc_hd__a21bo_2 _11479_ (.A1(_02389_),
    .A2(_02390_),
    .B1_N(_02416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02419_));
 sky130_fd_sc_hd__o211ai_2 _11480_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_02389_),
    .C1(_02390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02420_));
 sky130_fd_sc_hd__a22oi_2 _11481_ (.A1(_02308_),
    .A2(_02307_),
    .B1(_02271_),
    .B2(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02421_));
 sky130_fd_sc_hd__a21boi_2 _11482_ (.A1(_02270_),
    .A2(_02309_),
    .B1_N(_02310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02422_));
 sky130_fd_sc_hd__nand3_2 _11483_ (.A(_02419_),
    .B(_02420_),
    .C(_02422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02423_));
 sky130_fd_sc_hd__nand3_2 _11484_ (.A(_02417_),
    .B(_02421_),
    .C(_02418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02424_));
 sky130_fd_sc_hd__a21bo_2 _11485_ (.A1(_02423_),
    .A2(_02424_),
    .B1_N(_02354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02425_));
 sky130_fd_sc_hd__o211ai_2 _11486_ (.A1(_02351_),
    .A2(_02353_),
    .B1(_02423_),
    .C1(_02424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02426_));
 sky130_fd_sc_hd__nand2_2 _11487_ (.A(_02424_),
    .B(_02354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02427_));
 sky130_fd_sc_hd__nand3_2 _11488_ (.A(_02423_),
    .B(_02424_),
    .C(_02354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02428_));
 sky130_fd_sc_hd__a21o_2 _11489_ (.A1(_02423_),
    .A2(_02424_),
    .B1(_02354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02429_));
 sky130_fd_sc_hd__nand3_2 _11490_ (.A(_02429_),
    .B(_02336_),
    .C(_02428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02430_));
 sky130_fd_sc_hd__a21oi_2 _11491_ (.A1(_02428_),
    .A2(_02429_),
    .B1(_02336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02431_));
 sky130_fd_sc_hd__nand3_2 _11492_ (.A(_02337_),
    .B(_02425_),
    .C(_02426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02432_));
 sky130_fd_sc_hd__o2bb2ai_2 _11493_ (.A1_N(_02430_),
    .A2_N(_02432_),
    .B1(_02244_),
    .B2(_02245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02433_));
 sky130_fd_sc_hd__nand3b_2 _11494_ (.A_N(_02247_),
    .B(_02430_),
    .C(_02432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02434_));
 sky130_fd_sc_hd__nand2_2 _11495_ (.A(_02433_),
    .B(_02434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02435_));
 sky130_fd_sc_hd__a21o_2 _11496_ (.A1(_02323_),
    .A2(_02223_),
    .B1(_02321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02436_));
 sky130_fd_sc_hd__a21oi_2 _11497_ (.A1(_02323_),
    .A2(_02223_),
    .B1(_02321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02437_));
 sky130_fd_sc_hd__a21oi_2 _11498_ (.A1(_02433_),
    .A2(_02434_),
    .B1(_02436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02438_));
 sky130_fd_sc_hd__and3_2 _11499_ (.A(_02436_),
    .B(_02434_),
    .C(_02433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02439_));
 sky130_fd_sc_hd__nand3_2 _11500_ (.A(_02436_),
    .B(_02434_),
    .C(_02433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02440_));
 sky130_fd_sc_hd__o22ai_2 _11501_ (.A1(_02231_),
    .A2(_02328_),
    .B1(_02438_),
    .B2(_02439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02441_));
 sky130_fd_sc_hd__o31ai_2 _11502_ (.A1(_02231_),
    .A2(_02328_),
    .A3(_02438_),
    .B1(_02441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02442_));
 sky130_fd_sc_hd__o32a_2 _11503_ (.A1(_02141_),
    .A2(_02233_),
    .A3(_02328_),
    .B1(_02332_),
    .B2(_02334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02443_));
 sky130_fd_sc_hd__a21oi_2 _11504_ (.A1(_02442_),
    .A2(_02443_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02444_));
 sky130_fd_sc_hd__o21a_2 _11505_ (.A1(_02442_),
    .A2(_02443_),
    .B1(_02444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00285_));
 sky130_fd_sc_hd__o31a_2 _11506_ (.A1(_02242_),
    .A2(_02243_),
    .A3(_02245_),
    .B1(_02430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02445_));
 sky130_fd_sc_hd__o21ai_2 _11507_ (.A1(_02247_),
    .A2(_02431_),
    .B1(_02430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_2 _11508_ (.A(_02423_),
    .B(_02427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02447_));
 sky130_fd_sc_hd__a21boi_2 _11509_ (.A1(_02354_),
    .A2(_02424_),
    .B1_N(_02423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02448_));
 sky130_fd_sc_hd__o21ai_2 _11510_ (.A1(_02342_),
    .A2(_02341_),
    .B1(_02340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02449_));
 sky130_fd_sc_hd__o32a_2 _11511_ (.A1(_09624_),
    .A2(_09635_),
    .A3(_01860_),
    .B1(_02341_),
    .B2(_02342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02450_));
 sky130_fd_sc_hd__and2_2 _11512_ (.A(\a_h[1] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02451_));
 sky130_fd_sc_hd__nand2_2 _11513_ (.A(\a_h[1] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_2 _11514_ (.A(\a_h[2] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_2 _11515_ (.A(\a_h[3] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02454_));
 sky130_fd_sc_hd__nand4_2 _11516_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2_2 _11517_ (.A(_02453_),
    .B(_02454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02456_));
 sky130_fd_sc_hd__o211ai_2 _11518_ (.A1(_01871_),
    .A2(_02338_),
    .B1(_02452_),
    .C1(_02456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02457_));
 sky130_fd_sc_hd__a21o_2 _11519_ (.A1(_02455_),
    .A2(_02456_),
    .B1(_02452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02458_));
 sky130_fd_sc_hd__a22o_2 _11520_ (.A1(\a_h[1] ),
    .A2(\b_h[11] ),
    .B1(_02455_),
    .B2(_02456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02459_));
 sky130_fd_sc_hd__o2111ai_2 _11521_ (.A1(_01871_),
    .A2(_02338_),
    .B1(\a_h[1] ),
    .C1(\b_h[11] ),
    .D1(_02456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02460_));
 sky130_fd_sc_hd__nand3_2 _11522_ (.A(_02459_),
    .B(_02460_),
    .C(_02449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02461_));
 sky130_fd_sc_hd__and3_2 _11523_ (.A(_02450_),
    .B(_02457_),
    .C(_02458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02462_));
 sky130_fd_sc_hd__nand3_2 _11524_ (.A(_02450_),
    .B(_02457_),
    .C(_02458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02463_));
 sky130_fd_sc_hd__o2bb2ai_2 _11525_ (.A1_N(_02461_),
    .A2_N(_02463_),
    .B1(_09177_),
    .B2(_09657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02464_));
 sky130_fd_sc_hd__nand4_2 _11526_ (.A(_02463_),
    .B(\a_h[0] ),
    .C(_02461_),
    .D(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02465_));
 sky130_fd_sc_hd__o21ai_2 _11527_ (.A1(_02392_),
    .A2(_02406_),
    .B1(_02412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02466_));
 sky130_fd_sc_hd__a21oi_2 _11528_ (.A1(_02464_),
    .A2(_02465_),
    .B1(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02467_));
 sky130_fd_sc_hd__a21o_2 _11529_ (.A1(_02464_),
    .A2(_02465_),
    .B1(_02466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02468_));
 sky130_fd_sc_hd__and3_2 _11530_ (.A(_02464_),
    .B(_02466_),
    .C(_02465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02469_));
 sky130_fd_sc_hd__nand3_2 _11531_ (.A(_02464_),
    .B(_02466_),
    .C(_02465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02470_));
 sky130_fd_sc_hd__o21ai_2 _11532_ (.A1(_02467_),
    .A2(_02469_),
    .B1(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02471_));
 sky130_fd_sc_hd__nand4_2 _11533_ (.A(_02468_),
    .B(_02470_),
    .C(_02243_),
    .D(_02345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02472_));
 sky130_fd_sc_hd__o21bai_2 _11534_ (.A1(_02467_),
    .A2(_02469_),
    .B1_N(_02347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02473_));
 sky130_fd_sc_hd__nand3_2 _11535_ (.A(_02347_),
    .B(_02468_),
    .C(_02470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_2 _11536_ (.A(_02473_),
    .B(_02474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02475_));
 sky130_fd_sc_hd__nand2_2 _11537_ (.A(_02471_),
    .B(_02472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_2 _11538_ (.A(_02390_),
    .B(_02416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02477_));
 sky130_fd_sc_hd__a32oi_2 _11539_ (.A1(_02383_),
    .A2(_02384_),
    .A3(_02388_),
    .B1(_02390_),
    .B2(_02416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02478_));
 sky130_fd_sc_hd__nand2_2 _11540_ (.A(_02389_),
    .B(_02477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02479_));
 sky130_fd_sc_hd__a32oi_2 _11541_ (.A1(_02366_),
    .A2(_02368_),
    .A3(_02355_),
    .B1(_02379_),
    .B2(_02381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02480_));
 sky130_fd_sc_hd__o22ai_2 _11542_ (.A1(_02367_),
    .A2(_02371_),
    .B1(_02382_),
    .B2(_02369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02481_));
 sky130_fd_sc_hd__nor2_2 _11543_ (.A(_09449_),
    .B(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02482_));
 sky130_fd_sc_hd__a22oi_2 _11544_ (.A1(\a_h[9] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02483_));
 sky130_fd_sc_hd__a22o_2 _11545_ (.A1(\a_h[9] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02484_));
 sky130_fd_sc_hd__and4_2 _11546_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02485_));
 sky130_fd_sc_hd__nand4_2 _11547_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02486_));
 sky130_fd_sc_hd__o22ai_2 _11548_ (.A1(_09449_),
    .A2(_09602_),
    .B1(_02483_),
    .B2(_02485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02487_));
 sky130_fd_sc_hd__nand4_2 _11549_ (.A(_02484_),
    .B(_02486_),
    .C(\a_h[7] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02488_));
 sky130_fd_sc_hd__o21ai_2 _11550_ (.A1(_09449_),
    .A2(_09602_),
    .B1(_02486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02489_));
 sky130_fd_sc_hd__o21ai_2 _11551_ (.A1(_02483_),
    .A2(_02485_),
    .B1(_02482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02490_));
 sky130_fd_sc_hd__o21ai_2 _11552_ (.A1(_02483_),
    .A2(_02489_),
    .B1(_02490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_2 _11553_ (.A(_02487_),
    .B(_02488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02492_));
 sky130_fd_sc_hd__nand2_2 _11554_ (.A(_02357_),
    .B(_02364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02493_));
 sky130_fd_sc_hd__nand2_2 _11555_ (.A(_02361_),
    .B(_02493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02494_));
 sky130_fd_sc_hd__a21oi_2 _11556_ (.A1(_02357_),
    .A2(_02364_),
    .B1(_02360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02495_));
 sky130_fd_sc_hd__and2_2 _11557_ (.A(\a_h[10] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02496_));
 sky130_fd_sc_hd__nand2_2 _11558_ (.A(\a_h[10] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02497_));
 sky130_fd_sc_hd__nand2_2 _11559_ (.A(\a_h[11] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02498_));
 sky130_fd_sc_hd__nand2_2 _11560_ (.A(\a_h[12] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02499_));
 sky130_fd_sc_hd__a22oi_2 _11561_ (.A1(\a_h[12] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02500_));
 sky130_fd_sc_hd__nand2_2 _11562_ (.A(_02498_),
    .B(_02499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_2 _11563_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02502_));
 sky130_fd_sc_hd__nand4_2 _11564_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_2 _11565_ (.A(_02501_),
    .B(_02503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02504_));
 sky130_fd_sc_hd__nand2_2 _11566_ (.A(_02504_),
    .B(_02496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02505_));
 sky130_fd_sc_hd__o311a_2 _11567_ (.A1(_09526_),
    .A2(_09581_),
    .A3(_02502_),
    .B1(_02501_),
    .C1(_02497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02506_));
 sky130_fd_sc_hd__o211ai_2 _11568_ (.A1(_09482_),
    .A2(_09592_),
    .B1(_02501_),
    .C1(_02503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02507_));
 sky130_fd_sc_hd__o2bb2ai_2 _11569_ (.A1_N(_02501_),
    .A2_N(_02503_),
    .B1(_09482_),
    .B2(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02508_));
 sky130_fd_sc_hd__o21ai_2 _11570_ (.A1(_02498_),
    .A2(_02499_),
    .B1(_02496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02509_));
 sky130_fd_sc_hd__o211ai_2 _11571_ (.A1(_02509_),
    .A2(_02500_),
    .B1(_02495_),
    .C1(_02508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02510_));
 sky130_fd_sc_hd__a31o_2 _11572_ (.A1(_02504_),
    .A2(\b_h[2] ),
    .A3(\a_h[10] ),
    .B1(_02495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02511_));
 sky130_fd_sc_hd__nand3_2 _11573_ (.A(_02505_),
    .B(_02507_),
    .C(_02494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02512_));
 sky130_fd_sc_hd__nand2_2 _11574_ (.A(_02510_),
    .B(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02513_));
 sky130_fd_sc_hd__o2111ai_2 _11575_ (.A1(_02483_),
    .A2(_02489_),
    .B1(_02490_),
    .C1(_02510_),
    .D1(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_2 _11576_ (.A(_02513_),
    .B(_02491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02515_));
 sky130_fd_sc_hd__nand4_2 _11577_ (.A(_02487_),
    .B(_02488_),
    .C(_02510_),
    .D(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02516_));
 sky130_fd_sc_hd__o211a_2 _11578_ (.A1(_02483_),
    .A2(_02489_),
    .B1(_02490_),
    .C1(_02513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02517_));
 sky130_fd_sc_hd__a22o_2 _11579_ (.A1(_02487_),
    .A2(_02488_),
    .B1(_02510_),
    .B2(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02518_));
 sky130_fd_sc_hd__o211ai_2 _11580_ (.A1(_02369_),
    .A2(_02480_),
    .B1(_02514_),
    .C1(_02515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_2 _11581_ (.A(_02481_),
    .B(_02516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02520_));
 sky130_fd_sc_hd__nand3_2 _11582_ (.A(_02518_),
    .B(_02481_),
    .C(_02516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02521_));
 sky130_fd_sc_hd__nand2_2 _11583_ (.A(\a_h[6] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02522_));
 sky130_fd_sc_hd__nand2_2 _11584_ (.A(_02397_),
    .B(_02522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_2 _11585_ (.A(\a_h[6] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02524_));
 sky130_fd_sc_hd__nand4_2 _11586_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02525_));
 sky130_fd_sc_hd__nand3_2 _11587_ (.A(_02522_),
    .B(\b_h[7] ),
    .C(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02526_));
 sky130_fd_sc_hd__nand3_2 _11588_ (.A(_02397_),
    .B(\b_h[6] ),
    .C(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02527_));
 sky130_fd_sc_hd__o211ai_2 _11589_ (.A1(_09417_),
    .A2(_09613_),
    .B1(_02526_),
    .C1(_02527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02528_));
 sky130_fd_sc_hd__nand4_2 _11590_ (.A(_02523_),
    .B(_02525_),
    .C(\a_h[4] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02529_));
 sky130_fd_sc_hd__a21oi_2 _11591_ (.A1(_02373_),
    .A2(_02377_),
    .B1(_02375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02530_));
 sky130_fd_sc_hd__a21oi_2 _11592_ (.A1(_02528_),
    .A2(_02529_),
    .B1(_02530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02531_));
 sky130_fd_sc_hd__a21o_2 _11593_ (.A1(_02528_),
    .A2(_02529_),
    .B1(_02530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02532_));
 sky130_fd_sc_hd__nand3_2 _11594_ (.A(_02528_),
    .B(_02529_),
    .C(_02530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02533_));
 sky130_fd_sc_hd__and3_2 _11595_ (.A(_02396_),
    .B(\b_h[8] ),
    .C(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02534_));
 sky130_fd_sc_hd__a21oi_2 _11596_ (.A1(_02393_),
    .A2(_02396_),
    .B1(_02398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_2 _11597_ (.A1(_02532_),
    .A2(_02533_),
    .B1(_02535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02536_));
 sky130_fd_sc_hd__o2bb2ai_2 _11598_ (.A1_N(_02532_),
    .A2_N(_02533_),
    .B1(_02534_),
    .B2(_02398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02537_));
 sky130_fd_sc_hd__and3_2 _11599_ (.A(_02532_),
    .B(_02533_),
    .C(_02535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02538_));
 sky130_fd_sc_hd__nand4_2 _11600_ (.A(_02399_),
    .B(_02402_),
    .C(_02532_),
    .D(_02533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02539_));
 sky130_fd_sc_hd__nand2_2 _11601_ (.A(_02537_),
    .B(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02540_));
 sky130_fd_sc_hd__a21o_2 _11602_ (.A1(_02519_),
    .A2(_02521_),
    .B1(_02540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02541_));
 sky130_fd_sc_hd__o211ai_2 _11603_ (.A1(_02536_),
    .A2(_02538_),
    .B1(_02519_),
    .C1(_02521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02542_));
 sky130_fd_sc_hd__nand4_2 _11604_ (.A(_02519_),
    .B(_02521_),
    .C(_02537_),
    .D(_02539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02543_));
 sky130_fd_sc_hd__o2bb2ai_2 _11605_ (.A1_N(_02519_),
    .A2_N(_02521_),
    .B1(_02536_),
    .B2(_02538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02544_));
 sky130_fd_sc_hd__a21oi_2 _11606_ (.A1(_02543_),
    .A2(_02544_),
    .B1(_02479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02545_));
 sky130_fd_sc_hd__nand3_2 _11607_ (.A(_02541_),
    .B(_02542_),
    .C(_02478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02546_));
 sky130_fd_sc_hd__nand3_2 _11608_ (.A(_02479_),
    .B(_02543_),
    .C(_02544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02547_));
 sky130_fd_sc_hd__a21o_2 _11609_ (.A1(_02546_),
    .A2(_02547_),
    .B1(_02476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02548_));
 sky130_fd_sc_hd__nand4_2 _11610_ (.A(_02473_),
    .B(_02474_),
    .C(_02546_),
    .D(_02547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_2 _11611_ (.A(_02475_),
    .B(_02547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02550_));
 sky130_fd_sc_hd__a22o_2 _11612_ (.A1(_02471_),
    .A2(_02472_),
    .B1(_02546_),
    .B2(_02547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02551_));
 sky130_fd_sc_hd__a21oi_2 _11613_ (.A1(_02548_),
    .A2(_02549_),
    .B1(_02448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02552_));
 sky130_fd_sc_hd__o211ai_2 _11614_ (.A1(_02545_),
    .A2(_02550_),
    .B1(_02447_),
    .C1(_02551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02553_));
 sky130_fd_sc_hd__nand3_2 _11615_ (.A(_02448_),
    .B(_02548_),
    .C(_02549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02554_));
 sky130_fd_sc_hd__o2bb2ai_2 _11616_ (.A1_N(_02553_),
    .A2_N(_02554_),
    .B1(_02348_),
    .B2(_02350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02555_));
 sky130_fd_sc_hd__a31oi_2 _11617_ (.A1(_02448_),
    .A2(_02548_),
    .A3(_02549_),
    .B1(_02352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02556_));
 sky130_fd_sc_hd__nand3_2 _11618_ (.A(_02553_),
    .B(_02554_),
    .C(_02351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02557_));
 sky130_fd_sc_hd__a21o_2 _11619_ (.A1(_02553_),
    .A2(_02554_),
    .B1(_02352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02558_));
 sky130_fd_sc_hd__o211ai_2 _11620_ (.A1(_02348_),
    .A2(_02350_),
    .B1(_02553_),
    .C1(_02554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02559_));
 sky130_fd_sc_hd__nand3_2 _11621_ (.A(_02446_),
    .B(_02555_),
    .C(_02557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02560_));
 sky130_fd_sc_hd__a21oi_2 _11622_ (.A1(_02555_),
    .A2(_02557_),
    .B1(_02446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02561_));
 sky130_fd_sc_hd__o211ai_2 _11623_ (.A1(_02431_),
    .A2(_02445_),
    .B1(_02558_),
    .C1(_02559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02562_));
 sky130_fd_sc_hd__a2bb2oi_2 _11624_ (.A1_N(_02435_),
    .A2_N(_02437_),
    .B1(_02560_),
    .B2(_02562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_2 _11625_ (.A(_02440_),
    .B(_02561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02564_));
 sky130_fd_sc_hd__a21oi_2 _11626_ (.A1(_02564_),
    .A2(_02560_),
    .B1(_02563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02565_));
 sky130_fd_sc_hd__a21o_2 _11627_ (.A1(_02564_),
    .A2(_02560_),
    .B1(_02563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02566_));
 sky130_fd_sc_hd__o22ai_2 _11628_ (.A1(_02331_),
    .A2(_02438_),
    .B1(_02332_),
    .B2(_02334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_2 _11629_ (.A(_02441_),
    .B(_02567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02568_));
 sky130_fd_sc_hd__and3_2 _11630_ (.A(_02565_),
    .B(_02567_),
    .C(_02441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02569_));
 sky130_fd_sc_hd__a31o_2 _11631_ (.A1(_02565_),
    .A2(_02567_),
    .A3(_02441_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02570_));
 sky130_fd_sc_hd__a21oi_2 _11632_ (.A1(_02566_),
    .A2(_02568_),
    .B1(_02570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00286_));
 sky130_fd_sc_hd__a31o_2 _11633_ (.A1(_02439_),
    .A2(_02560_),
    .A3(_02562_),
    .B1(_02569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02571_));
 sky130_fd_sc_hd__a21oi_2 _11634_ (.A1(_02475_),
    .A2(_02547_),
    .B1(_02545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02572_));
 sky130_fd_sc_hd__a21o_2 _11635_ (.A1(_02475_),
    .A2(_02547_),
    .B1(_02545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02573_));
 sky130_fd_sc_hd__o31ai_2 _11636_ (.A1(_09177_),
    .A2(_09657_),
    .A3(_02462_),
    .B1(_02461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02574_));
 sky130_fd_sc_hd__o21ai_2 _11637_ (.A1(_02535_),
    .A2(_02531_),
    .B1(_02533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02575_));
 sky130_fd_sc_hd__o2bb2ai_2 _11638_ (.A1_N(_02451_),
    .A2_N(_02456_),
    .B1(_01871_),
    .B2(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02576_));
 sky130_fd_sc_hd__a21boi_2 _11639_ (.A1(_02456_),
    .A2(_02451_),
    .B1_N(_02455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_2 _11640_ (.A(\a_h[2] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02578_));
 sky130_fd_sc_hd__a22oi_2 _11641_ (.A1(\a_h[4] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02579_));
 sky130_fd_sc_hd__nor2_2 _11642_ (.A(_01888_),
    .B(_02338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02580_));
 sky130_fd_sc_hd__o21ai_2 _11643_ (.A1(_01888_),
    .A2(_02338_),
    .B1(_02578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02581_));
 sky130_fd_sc_hd__o21bai_2 _11644_ (.A1(_02579_),
    .A2(_02580_),
    .B1_N(_02578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02582_));
 sky130_fd_sc_hd__a41o_2 _11645_ (.A1(\a_h[3] ),
    .A2(\a_h[4] ),
    .A3(\b_h[9] ),
    .A4(\b_h[10] ),
    .B1(_02578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02583_));
 sky130_fd_sc_hd__o21ai_2 _11646_ (.A1(_02579_),
    .A2(_02580_),
    .B1(_02578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02584_));
 sky130_fd_sc_hd__o211ai_2 _11647_ (.A1(_02579_),
    .A2(_02583_),
    .B1(_02576_),
    .C1(_02584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02585_));
 sky130_fd_sc_hd__o211ai_2 _11648_ (.A1(_02581_),
    .A2(_02579_),
    .B1(_02577_),
    .C1(_02582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02586_));
 sky130_fd_sc_hd__nand2_2 _11649_ (.A(_02585_),
    .B(_02586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02587_));
 sky130_fd_sc_hd__and2_2 _11650_ (.A(\b_h[12] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02588_));
 sky130_fd_sc_hd__nand2_2 _11651_ (.A(\b_h[12] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02589_));
 sky130_fd_sc_hd__or2_2 _11652_ (.A(_01855_),
    .B(_02589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02590_));
 sky130_fd_sc_hd__a22oi_2 _11653_ (.A1(\a_h[1] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02591_));
 sky130_fd_sc_hd__a31oi_2 _11654_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_02588_),
    .B1(_02591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02592_));
 sky130_fd_sc_hd__a31o_2 _11655_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_02588_),
    .B1(_02591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_2 _11656_ (.A(_02587_),
    .B(_02592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02594_));
 sky130_fd_sc_hd__nand3_2 _11657_ (.A(_02585_),
    .B(_02586_),
    .C(_02593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02595_));
 sky130_fd_sc_hd__a21o_2 _11658_ (.A1(_02585_),
    .A2(_02586_),
    .B1(_02592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02596_));
 sky130_fd_sc_hd__nand3_2 _11659_ (.A(_02585_),
    .B(_02586_),
    .C(_02592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02597_));
 sky130_fd_sc_hd__a21oi_2 _11660_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02598_));
 sky130_fd_sc_hd__nand3b_2 _11661_ (.A_N(_02575_),
    .B(_02594_),
    .C(_02595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02599_));
 sky130_fd_sc_hd__nand3_2 _11662_ (.A(_02596_),
    .B(_02597_),
    .C(_02575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02600_));
 sky130_fd_sc_hd__nand2_2 _11663_ (.A(_02600_),
    .B(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02601_));
 sky130_fd_sc_hd__nand3_2 _11664_ (.A(_02599_),
    .B(_02600_),
    .C(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02602_));
 sky130_fd_sc_hd__a21o_2 _11665_ (.A1(_02599_),
    .A2(_02600_),
    .B1(_02574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02603_));
 sky130_fd_sc_hd__o21ai_2 _11666_ (.A1(_02598_),
    .A2(_02601_),
    .B1(_02603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02604_));
 sky130_fd_sc_hd__o2bb2ai_2 _11667_ (.A1_N(_02492_),
    .A2_N(_02510_),
    .B1(_02506_),
    .B2(_02511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02605_));
 sky130_fd_sc_hd__a21boi_2 _11668_ (.A1(_02492_),
    .A2(_02510_),
    .B1_N(_02512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02606_));
 sky130_fd_sc_hd__and2_2 _11669_ (.A(\a_h[11] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02607_));
 sky130_fd_sc_hd__nand2_2 _11670_ (.A(\a_h[11] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_2 _11671_ (.A(\a_h[12] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02609_));
 sky130_fd_sc_hd__nand2_2 _11672_ (.A(\a_h[13] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02610_));
 sky130_fd_sc_hd__a22oi_2 _11673_ (.A1(\a_h[13] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_2 _11674_ (.A(_02609_),
    .B(_02610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02612_));
 sky130_fd_sc_hd__nand2_2 _11675_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02613_));
 sky130_fd_sc_hd__nand4_2 _11676_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02614_));
 sky130_fd_sc_hd__nand2_2 _11677_ (.A(_02612_),
    .B(_02614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_2 _11678_ (.A(_02608_),
    .B(_02614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_2 _11679_ (.A(_02615_),
    .B(_02607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02617_));
 sky130_fd_sc_hd__a21o_2 _11680_ (.A1(_02612_),
    .A2(_02614_),
    .B1(_02607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02618_));
 sky130_fd_sc_hd__o2111ai_2 _11681_ (.A1(_01857_),
    .A2(_02613_),
    .B1(\a_h[11] ),
    .C1(\b_h[2] ),
    .D1(_02612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02619_));
 sky130_fd_sc_hd__a21o_2 _11682_ (.A1(_02497_),
    .A2(_02503_),
    .B1(_02500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02620_));
 sky130_fd_sc_hd__a21oi_2 _11683_ (.A1(_02497_),
    .A2(_02503_),
    .B1(_02500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02621_));
 sky130_fd_sc_hd__a21oi_2 _11684_ (.A1(_02618_),
    .A2(_02619_),
    .B1(_02621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02622_));
 sky130_fd_sc_hd__o211ai_2 _11685_ (.A1(_02611_),
    .A2(_02616_),
    .B1(_02620_),
    .C1(_02617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02623_));
 sky130_fd_sc_hd__nand3_2 _11686_ (.A(_02618_),
    .B(_02619_),
    .C(_02621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02624_));
 sky130_fd_sc_hd__nand2_2 _11687_ (.A(_02623_),
    .B(_02624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02625_));
 sky130_fd_sc_hd__nand2_2 _11688_ (.A(\a_h[8] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02626_));
 sky130_fd_sc_hd__a22oi_2 _11689_ (.A1(\a_h[10] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_2 _11690_ (.A(\a_h[10] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02628_));
 sky130_fd_sc_hd__and4_2 _11691_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02629_));
 sky130_fd_sc_hd__nand4_2 _11692_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02630_));
 sky130_fd_sc_hd__o22a_2 _11693_ (.A1(_09460_),
    .A2(_09602_),
    .B1(_02627_),
    .B2(_02629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02631_));
 sky130_fd_sc_hd__o21ai_2 _11694_ (.A1(_02627_),
    .A2(_02629_),
    .B1(_02626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02632_));
 sky130_fd_sc_hd__a41o_2 _11695_ (.A1(\a_h[9] ),
    .A2(\a_h[10] ),
    .A3(\b_h[3] ),
    .A4(\b_h[4] ),
    .B1(_02626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02633_));
 sky130_fd_sc_hd__and4b_2 _11696_ (.A_N(_02627_),
    .B(_02630_),
    .C(\a_h[8] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02634_));
 sky130_fd_sc_hd__o211ai_2 _11697_ (.A1(_02627_),
    .A2(_02629_),
    .B1(\a_h[8] ),
    .C1(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02635_));
 sky130_fd_sc_hd__o21ai_2 _11698_ (.A1(_09460_),
    .A2(_09602_),
    .B1(_02630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02636_));
 sky130_fd_sc_hd__o21ai_2 _11699_ (.A1(_02627_),
    .A2(_02636_),
    .B1(_02635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02637_));
 sky130_fd_sc_hd__o21ai_2 _11700_ (.A1(_02627_),
    .A2(_02633_),
    .B1(_02632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02638_));
 sky130_fd_sc_hd__o2111ai_2 _11701_ (.A1(_02627_),
    .A2(_02636_),
    .B1(_02635_),
    .C1(_02623_),
    .D1(_02624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02639_));
 sky130_fd_sc_hd__nand2_2 _11702_ (.A(_02625_),
    .B(_02637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02640_));
 sky130_fd_sc_hd__o2111ai_2 _11703_ (.A1(_02627_),
    .A2(_02633_),
    .B1(_02632_),
    .C1(_02623_),
    .D1(_02624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02641_));
 sky130_fd_sc_hd__inv_2 _11704_ (.A(_02641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02642_));
 sky130_fd_sc_hd__o2bb2ai_2 _11705_ (.A1_N(_02623_),
    .A2_N(_02624_),
    .B1(_02631_),
    .B2(_02634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02643_));
 sky130_fd_sc_hd__nand3_2 _11706_ (.A(_02640_),
    .B(_02605_),
    .C(_02639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02644_));
 sky130_fd_sc_hd__nand2_2 _11707_ (.A(_02606_),
    .B(_02643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02645_));
 sky130_fd_sc_hd__a21oi_2 _11708_ (.A1(_02639_),
    .A2(_02640_),
    .B1(_02605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02646_));
 sky130_fd_sc_hd__nand3_2 _11709_ (.A(_02606_),
    .B(_02641_),
    .C(_02643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02647_));
 sky130_fd_sc_hd__o21a_2 _11710_ (.A1(_02395_),
    .A2(_02524_),
    .B1(_02529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02648_));
 sky130_fd_sc_hd__nand2_2 _11711_ (.A(\a_h[7] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02649_));
 sky130_fd_sc_hd__nand2_2 _11712_ (.A(\a_h[7] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02650_));
 sky130_fd_sc_hd__nand4_2 _11713_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02651_));
 sky130_fd_sc_hd__nand2_2 _11714_ (.A(_02524_),
    .B(_02650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02652_));
 sky130_fd_sc_hd__nand3_2 _11715_ (.A(_02650_),
    .B(\b_h[7] ),
    .C(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02653_));
 sky130_fd_sc_hd__nand3_2 _11716_ (.A(_02524_),
    .B(\b_h[6] ),
    .C(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02654_));
 sky130_fd_sc_hd__nand4_2 _11717_ (.A(_02652_),
    .B(\b_h[8] ),
    .C(\a_h[5] ),
    .D(_02651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02655_));
 sky130_fd_sc_hd__o211ai_2 _11718_ (.A1(_09428_),
    .A2(_09613_),
    .B1(_02653_),
    .C1(_02654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02656_));
 sky130_fd_sc_hd__a22oi_2 _11719_ (.A1(_02484_),
    .A2(_02489_),
    .B1(_02655_),
    .B2(_02656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02657_));
 sky130_fd_sc_hd__o2111a_2 _11720_ (.A1(_02482_),
    .A2(_02485_),
    .B1(_02655_),
    .C1(_02656_),
    .D1(_02484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02658_));
 sky130_fd_sc_hd__o2111ai_2 _11721_ (.A1(_02482_),
    .A2(_02485_),
    .B1(_02655_),
    .C1(_02656_),
    .D1(_02484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02659_));
 sky130_fd_sc_hd__a211oi_2 _11722_ (.A1(_02525_),
    .A2(_02529_),
    .B1(_02657_),
    .C1(_02658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02660_));
 sky130_fd_sc_hd__o211a_2 _11723_ (.A1(_02657_),
    .A2(_02658_),
    .B1(_02525_),
    .C1(_02529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02661_));
 sky130_fd_sc_hd__o21bai_2 _11724_ (.A1(_02657_),
    .A2(_02658_),
    .B1_N(_02648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02662_));
 sky130_fd_sc_hd__nand3b_2 _11725_ (.A_N(_02657_),
    .B(_02659_),
    .C(_02648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02663_));
 sky130_fd_sc_hd__nand2_2 _11726_ (.A(_02662_),
    .B(_02663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02664_));
 sky130_fd_sc_hd__o2bb2ai_2 _11727_ (.A1_N(_02644_),
    .A2_N(_02647_),
    .B1(_02660_),
    .B2(_02661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_2 _11728_ (.A(_02644_),
    .B(_02664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02666_));
 sky130_fd_sc_hd__nand3_2 _11729_ (.A(_02644_),
    .B(_02647_),
    .C(_02664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02667_));
 sky130_fd_sc_hd__o2bb2ai_2 _11730_ (.A1_N(_02540_),
    .A2_N(_02519_),
    .B1(_02517_),
    .B2(_02520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02668_));
 sky130_fd_sc_hd__a21oi_2 _11731_ (.A1(_02665_),
    .A2(_02667_),
    .B1(_02668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02669_));
 sky130_fd_sc_hd__a21o_2 _11732_ (.A1(_02665_),
    .A2(_02667_),
    .B1(_02668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02670_));
 sky130_fd_sc_hd__o211a_2 _11733_ (.A1(_02646_),
    .A2(_02666_),
    .B1(_02668_),
    .C1(_02665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02671_));
 sky130_fd_sc_hd__o211ai_2 _11734_ (.A1(_02646_),
    .A2(_02666_),
    .B1(_02668_),
    .C1(_02665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02672_));
 sky130_fd_sc_hd__nand3_2 _11735_ (.A(_02604_),
    .B(_02670_),
    .C(_02672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02673_));
 sky130_fd_sc_hd__o21bai_2 _11736_ (.A1(_02669_),
    .A2(_02671_),
    .B1_N(_02604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02674_));
 sky130_fd_sc_hd__o21ai_2 _11737_ (.A1(_02669_),
    .A2(_02671_),
    .B1(_02604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02675_));
 sky130_fd_sc_hd__nand3b_2 _11738_ (.A_N(_02604_),
    .B(_02670_),
    .C(_02672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02676_));
 sky130_fd_sc_hd__nand3_2 _11739_ (.A(_02674_),
    .B(_02572_),
    .C(_02673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02677_));
 sky130_fd_sc_hd__a21oi_2 _11740_ (.A1(_02673_),
    .A2(_02674_),
    .B1(_02572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02678_));
 sky130_fd_sc_hd__nand3_2 _11741_ (.A(_02573_),
    .B(_02675_),
    .C(_02676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02679_));
 sky130_fd_sc_hd__a21oi_2 _11742_ (.A1(_02243_),
    .A2(_02345_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02680_));
 sky130_fd_sc_hd__a31o_2 _11743_ (.A1(_02468_),
    .A2(_02345_),
    .A3(_02243_),
    .B1(_02469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02681_));
 sky130_fd_sc_hd__o2bb2ai_2 _11744_ (.A1_N(_02677_),
    .A2_N(_02679_),
    .B1(_02680_),
    .B2(_02467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_2 _11745_ (.A(_02677_),
    .B(_02681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02683_));
 sky130_fd_sc_hd__a21bo_2 _11746_ (.A1(_02677_),
    .A2(_02679_),
    .B1_N(_02681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02684_));
 sky130_fd_sc_hd__o2111ai_2 _11747_ (.A1(_02347_),
    .A2(_02467_),
    .B1(_02470_),
    .C1(_02677_),
    .D1(_02679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02685_));
 sky130_fd_sc_hd__a21oi_2 _11748_ (.A1(_02554_),
    .A2(_02351_),
    .B1(_02552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02686_));
 sky130_fd_sc_hd__nand3_2 _11749_ (.A(_02684_),
    .B(_02685_),
    .C(_02686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02687_));
 sky130_fd_sc_hd__o221ai_2 _11750_ (.A1(_02678_),
    .A2(_02683_),
    .B1(_02552_),
    .B2(_02556_),
    .C1(_02682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02688_));
 sky130_fd_sc_hd__a21o_2 _11751_ (.A1(_02687_),
    .A2(_02688_),
    .B1(_02560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02689_));
 sky130_fd_sc_hd__nand3_2 _11752_ (.A(_02560_),
    .B(_02687_),
    .C(_02688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02690_));
 sky130_fd_sc_hd__nand2_2 _11753_ (.A(_02689_),
    .B(_02690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02691_));
 sky130_fd_sc_hd__a21oi_2 _11754_ (.A1(_02571_),
    .A2(_02691_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02692_));
 sky130_fd_sc_hd__o21a_2 _11755_ (.A1(_02571_),
    .A2(_02691_),
    .B1(_02692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00287_));
 sky130_fd_sc_hd__nand2_2 _11756_ (.A(_02679_),
    .B(_02683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02693_));
 sky130_fd_sc_hd__o21a_2 _11757_ (.A1(_02598_),
    .A2(_02601_),
    .B1(_02600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02694_));
 sky130_fd_sc_hd__a21oi_2 _11758_ (.A1(_02600_),
    .A2(_02602_),
    .B1(_02590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02695_));
 sky130_fd_sc_hd__and3_2 _11759_ (.A(_02590_),
    .B(_02600_),
    .C(_02602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02696_));
 sky130_fd_sc_hd__nor2_2 _11760_ (.A(_02695_),
    .B(_02696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02697_));
 sky130_fd_sc_hd__or2_2 _11761_ (.A(_02695_),
    .B(_02696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02698_));
 sky130_fd_sc_hd__a32oi_2 _11762_ (.A1(_02606_),
    .A2(_02641_),
    .A3(_02643_),
    .B1(_02644_),
    .B2(_02664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02699_));
 sky130_fd_sc_hd__o2bb2ai_2 _11763_ (.A1_N(_02664_),
    .A2_N(_02644_),
    .B1(_02642_),
    .B2(_02645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02700_));
 sky130_fd_sc_hd__o21a_2 _11764_ (.A1(_02524_),
    .A2(_02650_),
    .B1(_02655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02701_));
 sky130_fd_sc_hd__a21o_2 _11765_ (.A1(_02626_),
    .A2(_02630_),
    .B1(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02702_));
 sky130_fd_sc_hd__a21oi_2 _11766_ (.A1(_02626_),
    .A2(_02630_),
    .B1(_02627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_2 _11767_ (.A(\a_h[6] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_2 _11768_ (.A(\a_h[8] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02705_));
 sky130_fd_sc_hd__nand2_2 _11769_ (.A(_02649_),
    .B(_02705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02706_));
 sky130_fd_sc_hd__nand2_2 _11770_ (.A(\a_h[8] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02707_));
 sky130_fd_sc_hd__and4_2 _11771_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02708_));
 sky130_fd_sc_hd__nand4_2 _11772_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02709_));
 sky130_fd_sc_hd__o2bb2ai_2 _11773_ (.A1_N(_02706_),
    .A2_N(_02709_),
    .B1(_09439_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02710_));
 sky130_fd_sc_hd__o2111ai_2 _11774_ (.A1(_02650_),
    .A2(_02707_),
    .B1(\a_h[6] ),
    .C1(\b_h[8] ),
    .D1(_02706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02711_));
 sky130_fd_sc_hd__o221ai_2 _11775_ (.A1(_09439_),
    .A2(_09613_),
    .B1(_02650_),
    .B2(_02707_),
    .C1(_02706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02712_));
 sky130_fd_sc_hd__a21o_2 _11776_ (.A1(_02706_),
    .A2(_02709_),
    .B1(_02704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02713_));
 sky130_fd_sc_hd__nand3_2 _11777_ (.A(_02703_),
    .B(_02710_),
    .C(_02711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02714_));
 sky130_fd_sc_hd__a21oi_2 _11778_ (.A1(_02710_),
    .A2(_02711_),
    .B1(_02703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02715_));
 sky130_fd_sc_hd__nand3_2 _11779_ (.A(_02713_),
    .B(_02702_),
    .C(_02712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02716_));
 sky130_fd_sc_hd__a22o_2 _11780_ (.A1(_02651_),
    .A2(_02655_),
    .B1(_02714_),
    .B2(_02716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02717_));
 sky130_fd_sc_hd__o2111ai_2 _11781_ (.A1(_02524_),
    .A2(_02650_),
    .B1(_02655_),
    .C1(_02714_),
    .D1(_02716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02718_));
 sky130_fd_sc_hd__nand2_2 _11782_ (.A(_02717_),
    .B(_02718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02719_));
 sky130_fd_sc_hd__a21oi_2 _11783_ (.A1(_02624_),
    .A2(_02638_),
    .B1(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02720_));
 sky130_fd_sc_hd__a21o_2 _11784_ (.A1(_02624_),
    .A2(_02638_),
    .B1(_02622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02721_));
 sky130_fd_sc_hd__nand2_2 _11785_ (.A(\a_h[11] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02722_));
 sky130_fd_sc_hd__a22oi_2 _11786_ (.A1(\a_h[11] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_2 _11787_ (.A(_02628_),
    .B(_02722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_2 _11788_ (.A(\a_h[11] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02725_));
 sky130_fd_sc_hd__nand4_2 _11789_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02726_));
 sky130_fd_sc_hd__nand2_2 _11790_ (.A(\a_h[9] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02727_));
 sky130_fd_sc_hd__a22o_2 _11791_ (.A1(\a_h[9] ),
    .A2(\b_h[5] ),
    .B1(_02724_),
    .B2(_02726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02728_));
 sky130_fd_sc_hd__nand4_2 _11792_ (.A(_02724_),
    .B(_02726_),
    .C(\a_h[9] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_2 _11793_ (.A(_02728_),
    .B(_02729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02730_));
 sky130_fd_sc_hd__o22ai_2 _11794_ (.A1(_01857_),
    .A2(_02613_),
    .B1(_02608_),
    .B2(_02611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02731_));
 sky130_fd_sc_hd__nand2_2 _11795_ (.A(_02612_),
    .B(_02616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_2 _11796_ (.A(\a_h[12] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02733_));
 sky130_fd_sc_hd__nand2_2 _11797_ (.A(\a_h[13] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02734_));
 sky130_fd_sc_hd__nand2_2 _11798_ (.A(\a_h[14] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02735_));
 sky130_fd_sc_hd__a22oi_2 _11799_ (.A1(\a_h[14] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_2 _11800_ (.A(_02734_),
    .B(_02735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02737_));
 sky130_fd_sc_hd__nand2_2 _11801_ (.A(\a_h[14] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02738_));
 sky130_fd_sc_hd__nand4_2 _11802_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02739_));
 sky130_fd_sc_hd__nand2_2 _11803_ (.A(_02733_),
    .B(_02739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02740_));
 sky130_fd_sc_hd__a21o_2 _11804_ (.A1(_02737_),
    .A2(_02739_),
    .B1(_02733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02741_));
 sky130_fd_sc_hd__o2bb2ai_2 _11805_ (.A1_N(_02737_),
    .A2_N(_02739_),
    .B1(_09504_),
    .B2(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02742_));
 sky130_fd_sc_hd__o2111ai_2 _11806_ (.A1(_02610_),
    .A2(_02738_),
    .B1(\a_h[12] ),
    .C1(\b_h[2] ),
    .D1(_02737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02743_));
 sky130_fd_sc_hd__o211a_2 _11807_ (.A1(_02740_),
    .A2(_02736_),
    .B1(_02732_),
    .C1(_02741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02744_));
 sky130_fd_sc_hd__o211ai_2 _11808_ (.A1(_02740_),
    .A2(_02736_),
    .B1(_02732_),
    .C1(_02741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02745_));
 sky130_fd_sc_hd__nand3_2 _11809_ (.A(_02742_),
    .B(_02743_),
    .C(_02731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_2 _11810_ (.A(_02745_),
    .B(_02746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02747_));
 sky130_fd_sc_hd__nand4_2 _11811_ (.A(_02728_),
    .B(_02729_),
    .C(_02745_),
    .D(_02746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02748_));
 sky130_fd_sc_hd__nand2_2 _11812_ (.A(_02747_),
    .B(_02730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02749_));
 sky130_fd_sc_hd__a21o_2 _11813_ (.A1(_02745_),
    .A2(_02746_),
    .B1(_02730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02750_));
 sky130_fd_sc_hd__nand3_2 _11814_ (.A(_02745_),
    .B(_02746_),
    .C(_02730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02751_));
 sky130_fd_sc_hd__nand3_2 _11815_ (.A(_02749_),
    .B(_02720_),
    .C(_02748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02752_));
 sky130_fd_sc_hd__nand3_2 _11816_ (.A(_02721_),
    .B(_02750_),
    .C(_02751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_2 _11817_ (.A(_02752_),
    .B(_02753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02754_));
 sky130_fd_sc_hd__a21oi_2 _11818_ (.A1(_02752_),
    .A2(_02753_),
    .B1(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02755_));
 sky130_fd_sc_hd__nand3_2 _11819_ (.A(_02753_),
    .B(_02719_),
    .C(_02752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02756_));
 sky130_fd_sc_hd__nand4_2 _11820_ (.A(_02717_),
    .B(_02718_),
    .C(_02752_),
    .D(_02753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_2 _11821_ (.A(_02754_),
    .B(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02758_));
 sky130_fd_sc_hd__nand3_2 _11822_ (.A(_02758_),
    .B(_02699_),
    .C(_02757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02759_));
 sky130_fd_sc_hd__nand2_2 _11823_ (.A(_02700_),
    .B(_02756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02760_));
 sky130_fd_sc_hd__o21ai_2 _11824_ (.A1(_02755_),
    .A2(_02760_),
    .B1(_02759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02761_));
 sky130_fd_sc_hd__o21ai_2 _11825_ (.A1(_02648_),
    .A2(_02657_),
    .B1(_02659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02762_));
 sky130_fd_sc_hd__a22o_2 _11826_ (.A1(\a_h[2] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02763_));
 sky130_fd_sc_hd__and3_2 _11827_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(_02588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02764_));
 sky130_fd_sc_hd__nand4_2 _11828_ (.A(\a_h[1] ),
    .B(\a_h[2] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02765_));
 sky130_fd_sc_hd__a22oi_2 _11829_ (.A1(\a_h[0] ),
    .A2(\b_h[14] ),
    .B1(_02763_),
    .B2(_02765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02766_));
 sky130_fd_sc_hd__and4_2 _11830_ (.A(_02763_),
    .B(_02765_),
    .C(\a_h[0] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02767_));
 sky130_fd_sc_hd__nor2_2 _11831_ (.A(_02766_),
    .B(_02767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02768_));
 sky130_fd_sc_hd__o22ai_2 _11832_ (.A1(_01888_),
    .A2(_02338_),
    .B1(_02578_),
    .B2(_02579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_2 _11833_ (.A(\a_h[3] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_2 _11834_ (.A(\a_h[4] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02771_));
 sky130_fd_sc_hd__nand2_2 _11835_ (.A(\a_h[5] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02772_));
 sky130_fd_sc_hd__nand2_2 _11836_ (.A(_02771_),
    .B(_02772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_2 _11837_ (.A(\a_h[5] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02774_));
 sky130_fd_sc_hd__nand4_2 _11838_ (.A(\a_h[4] ),
    .B(\a_h[5] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02775_));
 sky130_fd_sc_hd__nand4_2 _11839_ (.A(_02773_),
    .B(_02775_),
    .C(\a_h[3] ),
    .D(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02776_));
 sky130_fd_sc_hd__a22o_2 _11840_ (.A1(\a_h[3] ),
    .A2(\b_h[11] ),
    .B1(_02773_),
    .B2(_02775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02777_));
 sky130_fd_sc_hd__o211ai_2 _11841_ (.A1(_09406_),
    .A2(_09646_),
    .B1(_02773_),
    .C1(_02775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02778_));
 sky130_fd_sc_hd__a21o_2 _11842_ (.A1(_02773_),
    .A2(_02775_),
    .B1(_02770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02779_));
 sky130_fd_sc_hd__nand3_2 _11843_ (.A(_02777_),
    .B(_02769_),
    .C(_02776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02780_));
 sky130_fd_sc_hd__a21oi_2 _11844_ (.A1(_02776_),
    .A2(_02777_),
    .B1(_02769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02781_));
 sky130_fd_sc_hd__nand3b_2 _11845_ (.A_N(_02769_),
    .B(_02778_),
    .C(_02779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02782_));
 sky130_fd_sc_hd__nand2_2 _11846_ (.A(_02780_),
    .B(_02782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02783_));
 sky130_fd_sc_hd__nand3_2 _11847_ (.A(_02768_),
    .B(_02780_),
    .C(_02782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02784_));
 sky130_fd_sc_hd__a2bb2o_2 _11848_ (.A1_N(_02766_),
    .A2_N(_02767_),
    .B1(_02780_),
    .B2(_02782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02785_));
 sky130_fd_sc_hd__nand2_2 _11849_ (.A(_02783_),
    .B(_02768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02786_));
 sky130_fd_sc_hd__o211ai_2 _11850_ (.A1(_02766_),
    .A2(_02767_),
    .B1(_02780_),
    .C1(_02782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02787_));
 sky130_fd_sc_hd__nand3_2 _11851_ (.A(_02785_),
    .B(_02762_),
    .C(_02784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02788_));
 sky130_fd_sc_hd__nand3b_2 _11852_ (.A_N(_02762_),
    .B(_02786_),
    .C(_02787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02789_));
 sky130_fd_sc_hd__nand2_2 _11853_ (.A(_02788_),
    .B(_02789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02790_));
 sky130_fd_sc_hd__a21boi_2 _11854_ (.A1(_02586_),
    .A2(_02592_),
    .B1_N(_02585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02791_));
 sky130_fd_sc_hd__inv_2 _11855_ (.A(_02791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02792_));
 sky130_fd_sc_hd__nand2_2 _11856_ (.A(_02790_),
    .B(_02792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02793_));
 sky130_fd_sc_hd__nand3_2 _11857_ (.A(_02788_),
    .B(_02789_),
    .C(_02791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02794_));
 sky130_fd_sc_hd__and2_2 _11858_ (.A(_02793_),
    .B(_02794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02795_));
 sky130_fd_sc_hd__nand2_2 _11859_ (.A(_02793_),
    .B(_02794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_2 _11860_ (.A(_02761_),
    .B(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02797_));
 sky130_fd_sc_hd__o211ai_2 _11861_ (.A1(_02755_),
    .A2(_02760_),
    .B1(_02759_),
    .C1(_02795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_2 _11862_ (.A(_02761_),
    .B(_02795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02799_));
 sky130_fd_sc_hd__o211ai_2 _11863_ (.A1(_02755_),
    .A2(_02760_),
    .B1(_02796_),
    .C1(_02759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02800_));
 sky130_fd_sc_hd__o21ai_2 _11864_ (.A1(_02604_),
    .A2(_02669_),
    .B1(_02672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02801_));
 sky130_fd_sc_hd__o21a_2 _11865_ (.A1(_02604_),
    .A2(_02669_),
    .B1(_02672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02802_));
 sky130_fd_sc_hd__nand3_2 _11866_ (.A(_02797_),
    .B(_02798_),
    .C(_02802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02803_));
 sky130_fd_sc_hd__nand3_2 _11867_ (.A(_02799_),
    .B(_02801_),
    .C(_02800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02804_));
 sky130_fd_sc_hd__a2bb2o_2 _11868_ (.A1_N(_02695_),
    .A2_N(_02696_),
    .B1(_02803_),
    .B2(_02804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02805_));
 sky130_fd_sc_hd__nand3_2 _11869_ (.A(_02803_),
    .B(_02804_),
    .C(_02697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02806_));
 sky130_fd_sc_hd__and3_2 _11870_ (.A(_02698_),
    .B(_02803_),
    .C(_02804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02807_));
 sky130_fd_sc_hd__a21oi_2 _11871_ (.A1(_02803_),
    .A2(_02804_),
    .B1(_02698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02808_));
 sky130_fd_sc_hd__nand3_2 _11872_ (.A(_02805_),
    .B(_02806_),
    .C(_02693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02809_));
 sky130_fd_sc_hd__inv_2 _11873_ (.A(_02809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02810_));
 sky130_fd_sc_hd__o31ai_2 _11874_ (.A1(_02693_),
    .A2(_02807_),
    .A3(_02808_),
    .B1(_02809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02811_));
 sky130_fd_sc_hd__nor2_2 _11875_ (.A(_02688_),
    .B(_02811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02812_));
 sky130_fd_sc_hd__and2_2 _11876_ (.A(_02688_),
    .B(_02811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02813_));
 sky130_fd_sc_hd__nor2_2 _11877_ (.A(_02812_),
    .B(_02813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02814_));
 sky130_fd_sc_hd__o21ai_2 _11878_ (.A1(_02435_),
    .A2(_02437_),
    .B1(_02560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02815_));
 sky130_fd_sc_hd__and3_2 _11879_ (.A(_02562_),
    .B(_02687_),
    .C(_02688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02816_));
 sky130_fd_sc_hd__nand2_2 _11880_ (.A(_02816_),
    .B(_02815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02817_));
 sky130_fd_sc_hd__nand4_2 _11881_ (.A(_02565_),
    .B(_02567_),
    .C(_02691_),
    .D(_02441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02818_));
 sky130_fd_sc_hd__a22o_2 _11882_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02569_),
    .B2(_02691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02819_));
 sky130_fd_sc_hd__a21oi_2 _11883_ (.A1(_02819_),
    .A2(_02814_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02820_));
 sky130_fd_sc_hd__o21a_2 _11884_ (.A1(_02814_),
    .A2(_02819_),
    .B1(_02820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00288_));
 sky130_fd_sc_hd__a32oi_2 _11885_ (.A1(_02797_),
    .A2(_02798_),
    .A3(_02802_),
    .B1(_02804_),
    .B2(_02698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02821_));
 sky130_fd_sc_hd__a21boi_2 _11886_ (.A1(_02803_),
    .A2(_02697_),
    .B1_N(_02804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02822_));
 sky130_fd_sc_hd__o2bb2ai_2 _11887_ (.A1_N(_02759_),
    .A2_N(_02796_),
    .B1(_02760_),
    .B2(_02755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02823_));
 sky130_fd_sc_hd__a2bb2oi_2 _11888_ (.A1_N(_02760_),
    .A2_N(_02755_),
    .B1(_02759_),
    .B2(_02796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02824_));
 sky130_fd_sc_hd__o21ai_2 _11889_ (.A1(_02701_),
    .A2(_02715_),
    .B1(_02714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02825_));
 sky130_fd_sc_hd__o21a_2 _11890_ (.A1(_02701_),
    .A2(_02715_),
    .B1(_02714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02826_));
 sky130_fd_sc_hd__a22o_2 _11891_ (.A1(\a_h[3] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02827_));
 sky130_fd_sc_hd__nand4_2 _11892_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02828_));
 sky130_fd_sc_hd__and3_2 _11893_ (.A(_02828_),
    .B(\b_h[14] ),
    .C(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02829_));
 sky130_fd_sc_hd__a22oi_2 _11894_ (.A1(\a_h[1] ),
    .A2(\b_h[14] ),
    .B1(_02827_),
    .B2(_02828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02830_));
 sky130_fd_sc_hd__a21oi_2 _11895_ (.A1(_02827_),
    .A2(_02829_),
    .B1(_02830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02831_));
 sky130_fd_sc_hd__a22oi_2 _11896_ (.A1(_02771_),
    .A2(_02772_),
    .B1(_02775_),
    .B2(_02770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02832_));
 sky130_fd_sc_hd__nand2_2 _11897_ (.A(\a_h[6] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02833_));
 sky130_fd_sc_hd__a22oi_2 _11898_ (.A1(\a_h[6] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2_2 _11899_ (.A(_02774_),
    .B(_02833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02835_));
 sky130_fd_sc_hd__nand2_2 _11900_ (.A(\a_h[6] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02836_));
 sky130_fd_sc_hd__nand4_2 _11901_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02837_));
 sky130_fd_sc_hd__nand2_2 _11902_ (.A(\a_h[4] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02838_));
 sky130_fd_sc_hd__o2bb2ai_2 _11903_ (.A1_N(_02835_),
    .A2_N(_02837_),
    .B1(_09417_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02839_));
 sky130_fd_sc_hd__o2111ai_2 _11904_ (.A1(_02772_),
    .A2(_02836_),
    .B1(\a_h[4] ),
    .C1(\b_h[11] ),
    .D1(_02835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02840_));
 sky130_fd_sc_hd__a21o_2 _11905_ (.A1(_02835_),
    .A2(_02837_),
    .B1(_02838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02841_));
 sky130_fd_sc_hd__o221ai_2 _11906_ (.A1(_09417_),
    .A2(_09646_),
    .B1(_02772_),
    .B2(_02836_),
    .C1(_02835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02842_));
 sky130_fd_sc_hd__nand3b_2 _11907_ (.A_N(_02832_),
    .B(_02841_),
    .C(_02842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02843_));
 sky130_fd_sc_hd__and3_2 _11908_ (.A(_02832_),
    .B(_02839_),
    .C(_02840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02844_));
 sky130_fd_sc_hd__nand3_2 _11909_ (.A(_02832_),
    .B(_02839_),
    .C(_02840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_2 _11910_ (.A(_02843_),
    .B(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02846_));
 sky130_fd_sc_hd__nand3_2 _11911_ (.A(_02831_),
    .B(_02843_),
    .C(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02847_));
 sky130_fd_sc_hd__a21o_2 _11912_ (.A1(_02843_),
    .A2(_02845_),
    .B1(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02848_));
 sky130_fd_sc_hd__nand3b_2 _11913_ (.A_N(_02831_),
    .B(_02843_),
    .C(_02845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_2 _11914_ (.A(_02846_),
    .B(_02831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02850_));
 sky130_fd_sc_hd__nand3_2 _11915_ (.A(_02848_),
    .B(_02825_),
    .C(_02847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02851_));
 sky130_fd_sc_hd__nand3_2 _11916_ (.A(_02826_),
    .B(_02849_),
    .C(_02850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02852_));
 sky130_fd_sc_hd__o21a_2 _11917_ (.A1(_02766_),
    .A2(_02767_),
    .B1(_02780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02853_));
 sky130_fd_sc_hd__a21bo_2 _11918_ (.A1(_02768_),
    .A2(_02782_),
    .B1_N(_02780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02854_));
 sky130_fd_sc_hd__o2bb2ai_2 _11919_ (.A1_N(_02851_),
    .A2_N(_02852_),
    .B1(_02853_),
    .B2(_02781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02855_));
 sky130_fd_sc_hd__nand2_2 _11920_ (.A(_02852_),
    .B(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02856_));
 sky130_fd_sc_hd__nand3_2 _11921_ (.A(_02851_),
    .B(_02852_),
    .C(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02857_));
 sky130_fd_sc_hd__nand2_2 _11922_ (.A(_02855_),
    .B(_02857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02858_));
 sky130_fd_sc_hd__nand2_2 _11923_ (.A(_02753_),
    .B(_02719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_2 _11924_ (.A(_02752_),
    .B(_02859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02860_));
 sky130_fd_sc_hd__a21boi_2 _11925_ (.A1(_02753_),
    .A2(_02719_),
    .B1_N(_02752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02861_));
 sky130_fd_sc_hd__nand2_2 _11926_ (.A(\a_h[9] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_2 _11927_ (.A(_02707_),
    .B(_02862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_2 _11928_ (.A(\a_h[9] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02864_));
 sky130_fd_sc_hd__nand4_2 _11929_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02865_));
 sky130_fd_sc_hd__nand4_2 _11930_ (.A(_02863_),
    .B(_02865_),
    .C(\a_h[7] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02866_));
 sky130_fd_sc_hd__nand3_2 _11931_ (.A(_02862_),
    .B(\b_h[7] ),
    .C(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02867_));
 sky130_fd_sc_hd__nand3_2 _11932_ (.A(_02707_),
    .B(\b_h[6] ),
    .C(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02868_));
 sky130_fd_sc_hd__o211ai_2 _11933_ (.A1(_09449_),
    .A2(_09613_),
    .B1(_02867_),
    .C1(_02868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02869_));
 sky130_fd_sc_hd__o21a_2 _11934_ (.A1(_02628_),
    .A2(_02722_),
    .B1(_02727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02870_));
 sky130_fd_sc_hd__o21ai_2 _11935_ (.A1(_02727_),
    .A2(_02723_),
    .B1(_02726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02871_));
 sky130_fd_sc_hd__o2bb2ai_2 _11936_ (.A1_N(_02866_),
    .A2_N(_02869_),
    .B1(_02870_),
    .B2(_02723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02872_));
 sky130_fd_sc_hd__nand3_2 _11937_ (.A(_02871_),
    .B(_02869_),
    .C(_02866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02873_));
 sky130_fd_sc_hd__a21oi_2 _11938_ (.A1(_02649_),
    .A2(_02705_),
    .B1(_02704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02874_));
 sky130_fd_sc_hd__a41o_2 _11939_ (.A1(\a_h[7] ),
    .A2(\a_h[8] ),
    .A3(\b_h[6] ),
    .A4(\b_h[7] ),
    .B1(_02874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02875_));
 sky130_fd_sc_hd__a21oi_2 _11940_ (.A1(_02872_),
    .A2(_02873_),
    .B1(_02875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02876_));
 sky130_fd_sc_hd__a211o_2 _11941_ (.A1(_02872_),
    .A2(_02873_),
    .B1(_02874_),
    .C1(_02708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02877_));
 sky130_fd_sc_hd__o211a_2 _11942_ (.A1(_02708_),
    .A2(_02874_),
    .B1(_02873_),
    .C1(_02872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02878_));
 sky130_fd_sc_hd__o211ai_2 _11943_ (.A1(_02708_),
    .A2(_02874_),
    .B1(_02873_),
    .C1(_02872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02879_));
 sky130_fd_sc_hd__nor2_2 _11944_ (.A(_02876_),
    .B(_02878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02880_));
 sky130_fd_sc_hd__a32oi_2 _11945_ (.A1(_02742_),
    .A2(_02743_),
    .A3(_02731_),
    .B1(_02729_),
    .B2(_02728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02881_));
 sky130_fd_sc_hd__a21oi_2 _11946_ (.A1(_02730_),
    .A2(_02746_),
    .B1(_02744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02882_));
 sky130_fd_sc_hd__nand2_2 _11947_ (.A(\a_h[10] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_2 _11948_ (.A(\a_h[12] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02884_));
 sky130_fd_sc_hd__a22oi_2 _11949_ (.A1(\a_h[12] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_2 _11950_ (.A(_02725_),
    .B(_02884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_2 _11951_ (.A(\a_h[12] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02887_));
 sky130_fd_sc_hd__nand4_2 _11952_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02888_));
 sky130_fd_sc_hd__a21o_2 _11953_ (.A1(_02886_),
    .A2(_02888_),
    .B1(_02883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02889_));
 sky130_fd_sc_hd__nand2_2 _11954_ (.A(_02883_),
    .B(_02888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02890_));
 sky130_fd_sc_hd__o21ai_2 _11955_ (.A1(_02885_),
    .A2(_02890_),
    .B1(_02889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02891_));
 sky130_fd_sc_hd__o21ai_2 _11956_ (.A1(_02733_),
    .A2(_02736_),
    .B1(_02739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_2 _11957_ (.A(_02737_),
    .B(_02740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02893_));
 sky130_fd_sc_hd__nor2_2 _11958_ (.A(_09515_),
    .B(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_2 _11959_ (.A(\a_h[13] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_2 _11960_ (.A(\a_h[15] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02896_));
 sky130_fd_sc_hd__a22oi_2 _11961_ (.A1(\a_h[15] ),
    .A2(\b_h[0] ),
    .B1(\b_h[1] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02897_));
 sky130_fd_sc_hd__nand2_2 _11962_ (.A(_02738_),
    .B(_02896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_2 _11963_ (.A(\a_h[15] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02899_));
 sky130_fd_sc_hd__nand4_2 _11964_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[0] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02900_));
 sky130_fd_sc_hd__nand2_2 _11965_ (.A(_02898_),
    .B(_02900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02901_));
 sky130_fd_sc_hd__o2bb2ai_2 _11966_ (.A1_N(_02898_),
    .A2_N(_02900_),
    .B1(_09515_),
    .B2(_09592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02902_));
 sky130_fd_sc_hd__o2111ai_2 _11967_ (.A1(_02735_),
    .A2(_02899_),
    .B1(\a_h[13] ),
    .C1(\b_h[2] ),
    .D1(_02898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_2 _11968_ (.A(_02895_),
    .B(_02900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_2 _11969_ (.A(_02901_),
    .B(_02894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02905_));
 sky130_fd_sc_hd__o211ai_2 _11970_ (.A1(_02904_),
    .A2(_02897_),
    .B1(_02893_),
    .C1(_02905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02906_));
 sky130_fd_sc_hd__nand3_2 _11971_ (.A(_02902_),
    .B(_02903_),
    .C(_02892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02907_));
 sky130_fd_sc_hd__nand2_2 _11972_ (.A(_02906_),
    .B(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02908_));
 sky130_fd_sc_hd__o211ai_2 _11973_ (.A1(_02890_),
    .A2(_02885_),
    .B1(_02889_),
    .C1(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02909_));
 sky130_fd_sc_hd__o2111a_2 _11974_ (.A1(_02890_),
    .A2(_02885_),
    .B1(_02889_),
    .C1(_02906_),
    .D1(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02910_));
 sky130_fd_sc_hd__o2111ai_2 _11975_ (.A1(_02890_),
    .A2(_02885_),
    .B1(_02889_),
    .C1(_02906_),
    .D1(_02907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02911_));
 sky130_fd_sc_hd__nand2_2 _11976_ (.A(_02908_),
    .B(_02891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02912_));
 sky130_fd_sc_hd__nand3_2 _11977_ (.A(_02906_),
    .B(_02907_),
    .C(_02891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02913_));
 sky130_fd_sc_hd__a21o_2 _11978_ (.A1(_02906_),
    .A2(_02907_),
    .B1(_02891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02914_));
 sky130_fd_sc_hd__o2bb2ai_2 _11979_ (.A1_N(_02891_),
    .A2_N(_02908_),
    .B1(_02744_),
    .B2(_02881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02915_));
 sky130_fd_sc_hd__o211ai_2 _11980_ (.A1(_02744_),
    .A2(_02881_),
    .B1(_02911_),
    .C1(_02912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02916_));
 sky130_fd_sc_hd__nand3_2 _11981_ (.A(_02882_),
    .B(_02913_),
    .C(_02914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02917_));
 sky130_fd_sc_hd__inv_2 _11982_ (.A(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02918_));
 sky130_fd_sc_hd__o21ai_2 _11983_ (.A1(_02910_),
    .A2(_02915_),
    .B1(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02919_));
 sky130_fd_sc_hd__nand2_2 _11984_ (.A(_02919_),
    .B(_02880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02920_));
 sky130_fd_sc_hd__o21ai_2 _11985_ (.A1(_02876_),
    .A2(_02878_),
    .B1(_02916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02921_));
 sky130_fd_sc_hd__o211a_2 _11986_ (.A1(_02876_),
    .A2(_02878_),
    .B1(_02916_),
    .C1(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02922_));
 sky130_fd_sc_hd__o211ai_2 _11987_ (.A1(_02910_),
    .A2(_02915_),
    .B1(_02917_),
    .C1(_02880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02923_));
 sky130_fd_sc_hd__a22o_2 _11988_ (.A1(_02877_),
    .A2(_02879_),
    .B1(_02916_),
    .B2(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02924_));
 sky130_fd_sc_hd__nand3_2 _11989_ (.A(_02924_),
    .B(_02860_),
    .C(_02923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02925_));
 sky130_fd_sc_hd__inv_2 _11990_ (.A(_02925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_2 _11991_ (.A(_02861_),
    .B(_02920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02927_));
 sky130_fd_sc_hd__o211ai_2 _11992_ (.A1(_02921_),
    .A2(_02918_),
    .B1(_02861_),
    .C1(_02920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_2 _11993_ (.A(_02925_),
    .B(_02928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_2 _11994_ (.A(_02928_),
    .B(_02858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02930_));
 sky130_fd_sc_hd__a21o_2 _11995_ (.A1(_02925_),
    .A2(_02928_),
    .B1(_02858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02931_));
 sky130_fd_sc_hd__nand4_2 _11996_ (.A(_02855_),
    .B(_02857_),
    .C(_02925_),
    .D(_02928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02932_));
 sky130_fd_sc_hd__inv_2 _11997_ (.A(_02932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_2 _11998_ (.A(_02929_),
    .B(_02858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02934_));
 sky130_fd_sc_hd__a21o_2 _11999_ (.A1(_02858_),
    .A2(_02929_),
    .B1(_02824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02935_));
 sky130_fd_sc_hd__nand3_2 _12000_ (.A(_02934_),
    .B(_02823_),
    .C(_02932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02936_));
 sky130_fd_sc_hd__o211ai_2 _12001_ (.A1(_02930_),
    .A2(_02926_),
    .B1(_02824_),
    .C1(_02931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02937_));
 sky130_fd_sc_hd__a31o_2 _12002_ (.A1(\a_h[0] ),
    .A2(\b_h[14] ),
    .A3(_02763_),
    .B1(_02764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02938_));
 sky130_fd_sc_hd__nand2_2 _12003_ (.A(_02788_),
    .B(_02791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02939_));
 sky130_fd_sc_hd__o211a_2 _12004_ (.A1(_02764_),
    .A2(_02767_),
    .B1(_02789_),
    .C1(_02939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02940_));
 sky130_fd_sc_hd__a21oi_2 _12005_ (.A1(_02789_),
    .A2(_02939_),
    .B1(_02938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02941_));
 sky130_fd_sc_hd__a32o_2 _12006_ (.A1(_02789_),
    .A2(_02938_),
    .A3(_02939_),
    .B1(\b_h[15] ),
    .B2(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02942_));
 sky130_fd_sc_hd__nor2_2 _12007_ (.A(_02941_),
    .B(_02942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02943_));
 sky130_fd_sc_hd__o211a_2 _12008_ (.A1(_02940_),
    .A2(_02941_),
    .B1(\a_h[0] ),
    .C1(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02944_));
 sky130_fd_sc_hd__o211ai_2 _12009_ (.A1(_02940_),
    .A2(_02941_),
    .B1(\a_h[0] ),
    .C1(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02945_));
 sky130_fd_sc_hd__o21ai_2 _12010_ (.A1(_02941_),
    .A2(_02942_),
    .B1(_02945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02946_));
 sky130_fd_sc_hd__o2bb2ai_2 _12011_ (.A1_N(_02936_),
    .A2_N(_02937_),
    .B1(_02943_),
    .B2(_02944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02947_));
 sky130_fd_sc_hd__o2111ai_2 _12012_ (.A1(_02941_),
    .A2(_02942_),
    .B1(_02945_),
    .C1(_02937_),
    .D1(_02936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02948_));
 sky130_fd_sc_hd__a21oi_2 _12013_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02949_));
 sky130_fd_sc_hd__a21o_2 _12014_ (.A1(_02936_),
    .A2(_02937_),
    .B1(_02946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02950_));
 sky130_fd_sc_hd__o211ai_2 _12015_ (.A1(_02943_),
    .A2(_02944_),
    .B1(_02936_),
    .C1(_02937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02951_));
 sky130_fd_sc_hd__nand2_2 _12016_ (.A(_02821_),
    .B(_02951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02952_));
 sky130_fd_sc_hd__and3_2 _12017_ (.A(_02950_),
    .B(_02951_),
    .C(_02821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02953_));
 sky130_fd_sc_hd__a21o_2 _12018_ (.A1(_02947_),
    .A2(_02948_),
    .B1(_02822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02954_));
 sky130_fd_sc_hd__nand3_2 _12019_ (.A(_02822_),
    .B(_02947_),
    .C(_02948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02955_));
 sky130_fd_sc_hd__o21ai_2 _12020_ (.A1(_02949_),
    .A2(_02952_),
    .B1(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02956_));
 sky130_fd_sc_hd__nand2_2 _12021_ (.A(_02955_),
    .B(_02695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ai_2 _12022_ (.A1(_02590_),
    .A2(_02694_),
    .B1(_02956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02958_));
 sky130_fd_sc_hd__o211ai_2 _12023_ (.A1(_02953_),
    .A2(_02957_),
    .B1(_02810_),
    .C1(_02958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02959_));
 sky130_fd_sc_hd__o21ai_2 _12024_ (.A1(_02590_),
    .A2(_02694_),
    .B1(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02960_));
 sky130_fd_sc_hd__nand2_2 _12025_ (.A(_02956_),
    .B(_02695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02961_));
 sky130_fd_sc_hd__o211a_2 _12026_ (.A1(_02960_),
    .A2(_02953_),
    .B1(_02809_),
    .C1(_02961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02962_));
 sky130_fd_sc_hd__o211ai_2 _12027_ (.A1(_02960_),
    .A2(_02953_),
    .B1(_02809_),
    .C1(_02961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02963_));
 sky130_fd_sc_hd__and2_2 _12028_ (.A(_02959_),
    .B(_02963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02964_));
 sky130_fd_sc_hd__a21o_2 _12029_ (.A1(_02819_),
    .A2(_02814_),
    .B1(_02812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02965_));
 sky130_fd_sc_hd__a21oi_2 _12030_ (.A1(_02965_),
    .A2(_02964_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02966_));
 sky130_fd_sc_hd__o21a_2 _12031_ (.A1(_02964_),
    .A2(_02965_),
    .B1(_02966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00289_));
 sky130_fd_sc_hd__a21boi_2 _12032_ (.A1(_02937_),
    .A2(_02946_),
    .B1_N(_02936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02967_));
 sky130_fd_sc_hd__o2bb2ai_2 _12033_ (.A1_N(_02937_),
    .A2_N(_02946_),
    .B1(_02933_),
    .B2(_02935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02968_));
 sky130_fd_sc_hd__nand2_2 _12034_ (.A(_02916_),
    .B(_02880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02969_));
 sky130_fd_sc_hd__o21ai_2 _12035_ (.A1(_02876_),
    .A2(_02878_),
    .B1(_02917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2_2 _12036_ (.A(_02917_),
    .B(_02969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_2 _12037_ (.A(_02886_),
    .B(_02890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02972_));
 sky130_fd_sc_hd__a21oi_2 _12038_ (.A1(_02883_),
    .A2(_02888_),
    .B1(_02885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02973_));
 sky130_fd_sc_hd__nor2_2 _12039_ (.A(_09460_),
    .B(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02974_));
 sky130_fd_sc_hd__nand2_2 _12040_ (.A(\a_h[8] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02975_));
 sky130_fd_sc_hd__nand2_2 _12041_ (.A(\a_h[10] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_2 _12042_ (.A(_02864_),
    .B(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_2 _12043_ (.A(\a_h[10] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02978_));
 sky130_fd_sc_hd__nand4_2 _12044_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02979_));
 sky130_fd_sc_hd__o2bb2ai_2 _12045_ (.A1_N(_02864_),
    .A2_N(_02976_),
    .B1(_02978_),
    .B2(_02862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02980_));
 sky130_fd_sc_hd__o21ai_2 _12046_ (.A1(_09460_),
    .A2(_09613_),
    .B1(_02980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02981_));
 sky130_fd_sc_hd__o2111ai_2 _12047_ (.A1(_02862_),
    .A2(_02978_),
    .B1(\a_h[8] ),
    .C1(\b_h[8] ),
    .D1(_02977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02982_));
 sky130_fd_sc_hd__o221ai_2 _12048_ (.A1(_09460_),
    .A2(_09613_),
    .B1(_02862_),
    .B2(_02978_),
    .C1(_02977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_2 _12049_ (.A(_02980_),
    .B(_02974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02984_));
 sky130_fd_sc_hd__and3_2 _12050_ (.A(_02984_),
    .B(_02972_),
    .C(_02983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02985_));
 sky130_fd_sc_hd__nand3_2 _12051_ (.A(_02984_),
    .B(_02972_),
    .C(_02983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02986_));
 sky130_fd_sc_hd__a21oi_2 _12052_ (.A1(_02983_),
    .A2(_02984_),
    .B1(_02972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02987_));
 sky130_fd_sc_hd__nand3_2 _12053_ (.A(_02973_),
    .B(_02981_),
    .C(_02982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02988_));
 sky130_fd_sc_hd__o21a_2 _12054_ (.A1(_02707_),
    .A2(_02862_),
    .B1(_02866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02989_));
 sky130_fd_sc_hd__o21ai_2 _12055_ (.A1(_02707_),
    .A2(_02862_),
    .B1(_02866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02990_));
 sky130_fd_sc_hd__a21oi_2 _12056_ (.A1(_02986_),
    .A2(_02988_),
    .B1(_02989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02991_));
 sky130_fd_sc_hd__a22o_2 _12057_ (.A1(_02865_),
    .A2(_02866_),
    .B1(_02986_),
    .B2(_02988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02992_));
 sky130_fd_sc_hd__nand2_2 _12058_ (.A(_02986_),
    .B(_02989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02993_));
 sky130_fd_sc_hd__nor2_2 _12059_ (.A(_02987_),
    .B(_02993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02994_));
 sky130_fd_sc_hd__o21ai_2 _12060_ (.A1(_02987_),
    .A2(_02993_),
    .B1(_02992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02995_));
 sky130_fd_sc_hd__nand2_2 _12061_ (.A(\a_h[14] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_2 _12062_ (.A(_02899_),
    .B(_02996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02997_));
 sky130_fd_sc_hd__nand4_2 _12063_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[1] ),
    .D(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_02998_));
 sky130_fd_sc_hd__and2_2 _12064_ (.A(_02997_),
    .B(_02998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_02999_));
 sky130_fd_sc_hd__nand2_2 _12065_ (.A(_02997_),
    .B(_02998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03000_));
 sky130_fd_sc_hd__a21oi_2 _12066_ (.A1(_02895_),
    .A2(_02900_),
    .B1(_02897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03001_));
 sky130_fd_sc_hd__nand4_2 _12067_ (.A(_02898_),
    .B(_02904_),
    .C(_02997_),
    .D(_02998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03002_));
 sky130_fd_sc_hd__o211ai_2 _12068_ (.A1(_02895_),
    .A2(_02897_),
    .B1(_02900_),
    .C1(_03000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03003_));
 sky130_fd_sc_hd__inv_2 _12069_ (.A(_03003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_2 _12070_ (.A(_03002_),
    .B(_03003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03005_));
 sky130_fd_sc_hd__nand2_2 _12071_ (.A(\a_h[11] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_2 _12072_ (.A(\a_h[13] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_2 _12073_ (.A(\a_h[13] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03008_));
 sky130_fd_sc_hd__nand4_2 _12074_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03009_));
 sky130_fd_sc_hd__a22oi_2 _12075_ (.A1(\a_h[13] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_2 _12076_ (.A(_02887_),
    .B(_03008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03011_));
 sky130_fd_sc_hd__a22oi_2 _12077_ (.A1(\a_h[11] ),
    .A2(\b_h[5] ),
    .B1(_03009_),
    .B2(_03011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03012_));
 sky130_fd_sc_hd__a22o_2 _12078_ (.A1(\a_h[11] ),
    .A2(\b_h[5] ),
    .B1(_03009_),
    .B2(_03011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03013_));
 sky130_fd_sc_hd__and4_2 _12079_ (.A(_03011_),
    .B(\b_h[5] ),
    .C(\a_h[11] ),
    .D(_03009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03014_));
 sky130_fd_sc_hd__o2111ai_2 _12080_ (.A1(_02884_),
    .A2(_03007_),
    .B1(\a_h[11] ),
    .C1(\b_h[5] ),
    .D1(_03011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03015_));
 sky130_fd_sc_hd__o221ai_2 _12081_ (.A1(_09493_),
    .A2(_09602_),
    .B1(_02884_),
    .B2(_03007_),
    .C1(_03011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03016_));
 sky130_fd_sc_hd__a21o_2 _12082_ (.A1(_03009_),
    .A2(_03011_),
    .B1(_03006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_2 _12083_ (.A(_03016_),
    .B(_03017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03018_));
 sky130_fd_sc_hd__o2bb2ai_2 _12084_ (.A1_N(_03002_),
    .A2_N(_03003_),
    .B1(_03012_),
    .B2(_03014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03019_));
 sky130_fd_sc_hd__nand4_2 _12085_ (.A(_03002_),
    .B(_03003_),
    .C(_03013_),
    .D(_03015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03020_));
 sky130_fd_sc_hd__nand2_2 _12086_ (.A(_03005_),
    .B(_03018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03021_));
 sky130_fd_sc_hd__a22oi_2 _12087_ (.A1(_02999_),
    .A2(_03001_),
    .B1(_03013_),
    .B2(_03015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03022_));
 sky130_fd_sc_hd__o21ai_2 _12088_ (.A1(_03012_),
    .A2(_03014_),
    .B1(_03002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03023_));
 sky130_fd_sc_hd__nand4_2 _12089_ (.A(_03002_),
    .B(_03003_),
    .C(_03016_),
    .D(_03017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_2 _12090_ (.A(_02906_),
    .B(_02891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03025_));
 sky130_fd_sc_hd__nand4_2 _12091_ (.A(_02906_),
    .B(_02909_),
    .C(_03019_),
    .D(_03020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03026_));
 sky130_fd_sc_hd__nand4_2 _12092_ (.A(_02907_),
    .B(_03021_),
    .C(_03024_),
    .D(_03025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03027_));
 sky130_fd_sc_hd__o21ai_2 _12093_ (.A1(_02991_),
    .A2(_02994_),
    .B1(_03027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03028_));
 sky130_fd_sc_hd__o211a_2 _12094_ (.A1(_02991_),
    .A2(_02994_),
    .B1(_03026_),
    .C1(_03027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03029_));
 sky130_fd_sc_hd__o211ai_2 _12095_ (.A1(_02991_),
    .A2(_02994_),
    .B1(_03026_),
    .C1(_03027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03030_));
 sky130_fd_sc_hd__a21oi_2 _12096_ (.A1(_03026_),
    .A2(_03027_),
    .B1(_02995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03031_));
 sky130_fd_sc_hd__a21o_2 _12097_ (.A1(_03026_),
    .A2(_03027_),
    .B1(_02995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03032_));
 sky130_fd_sc_hd__nand2_2 _12098_ (.A(_03026_),
    .B(_03028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03033_));
 sky130_fd_sc_hd__a21oi_2 _12099_ (.A1(_03030_),
    .A2(_03032_),
    .B1(_02971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03034_));
 sky130_fd_sc_hd__o2bb2ai_2 _12100_ (.A1_N(_02916_),
    .A2_N(_02970_),
    .B1(_03029_),
    .B2(_03031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03035_));
 sky130_fd_sc_hd__a21oi_2 _12101_ (.A1(_02917_),
    .A2(_02969_),
    .B1(_03029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03036_));
 sky130_fd_sc_hd__nand3_2 _12102_ (.A(_02971_),
    .B(_03030_),
    .C(_03032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03037_));
 sky130_fd_sc_hd__a21bo_2 _12103_ (.A1(_02872_),
    .A2(_02875_),
    .B1_N(_02873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03038_));
 sky130_fd_sc_hd__a21boi_2 _12104_ (.A1(_02872_),
    .A2(_02875_),
    .B1_N(_02873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_2 _12105_ (.A(\a_h[3] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03040_));
 sky130_fd_sc_hd__nand2_2 _12106_ (.A(\a_h[4] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03041_));
 sky130_fd_sc_hd__nand2_2 _12107_ (.A(_03040_),
    .B(_03041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03042_));
 sky130_fd_sc_hd__nand2_2 _12108_ (.A(\a_h[4] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03043_));
 sky130_fd_sc_hd__nand4_2 _12109_ (.A(\a_h[3] ),
    .B(\a_h[4] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03044_));
 sky130_fd_sc_hd__and4_2 _12110_ (.A(_03042_),
    .B(_03044_),
    .C(\a_h[2] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03045_));
 sky130_fd_sc_hd__a22oi_2 _12111_ (.A1(\a_h[2] ),
    .A2(\b_h[14] ),
    .B1(_03042_),
    .B2(_03044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03046_));
 sky130_fd_sc_hd__nor2_2 _12112_ (.A(_03045_),
    .B(_03046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03047_));
 sky130_fd_sc_hd__a21o_2 _12113_ (.A1(_02837_),
    .A2(_02838_),
    .B1(_02834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03048_));
 sky130_fd_sc_hd__a21oi_2 _12114_ (.A1(_02837_),
    .A2(_02838_),
    .B1(_02834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_2 _12115_ (.A(\a_h[5] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_2 _12116_ (.A(\a_h[7] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03051_));
 sky130_fd_sc_hd__a22oi_2 _12117_ (.A1(\a_h[7] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2_2 _12118_ (.A(_02836_),
    .B(_03051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_2 _12119_ (.A(\a_h[7] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03054_));
 sky130_fd_sc_hd__nand4_2 _12120_ (.A(\a_h[6] ),
    .B(\a_h[7] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03055_));
 sky130_fd_sc_hd__o21ai_2 _12121_ (.A1(_02836_),
    .A2(_03051_),
    .B1(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03056_));
 sky130_fd_sc_hd__a21o_2 _12122_ (.A1(_03053_),
    .A2(_03055_),
    .B1(_03050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03057_));
 sky130_fd_sc_hd__o2bb2ai_2 _12123_ (.A1_N(_03053_),
    .A2_N(_03055_),
    .B1(_09428_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03058_));
 sky130_fd_sc_hd__nand3_2 _12124_ (.A(_03055_),
    .B(\b_h[11] ),
    .C(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03059_));
 sky130_fd_sc_hd__o211a_2 _12125_ (.A1(_03052_),
    .A2(_03056_),
    .B1(_03048_),
    .C1(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03060_));
 sky130_fd_sc_hd__o211ai_2 _12126_ (.A1(_03052_),
    .A2(_03056_),
    .B1(_03048_),
    .C1(_03057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03061_));
 sky130_fd_sc_hd__o211ai_2 _12127_ (.A1(_03059_),
    .A2(_03052_),
    .B1(_03049_),
    .C1(_03058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_2 _12128_ (.A(_03061_),
    .B(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03063_));
 sky130_fd_sc_hd__o21ai_2 _12129_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03064_));
 sky130_fd_sc_hd__nand3_2 _12130_ (.A(_03047_),
    .B(_03061_),
    .C(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03065_));
 sky130_fd_sc_hd__o21ai_2 _12131_ (.A1(_03045_),
    .A2(_03046_),
    .B1(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03066_));
 sky130_fd_sc_hd__nand2_2 _12132_ (.A(_03063_),
    .B(_03047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03067_));
 sky130_fd_sc_hd__nand3_2 _12133_ (.A(_03038_),
    .B(_03064_),
    .C(_03065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03068_));
 sky130_fd_sc_hd__o211ai_2 _12134_ (.A1(_03066_),
    .A2(_03060_),
    .B1(_03039_),
    .C1(_03067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_2 _12135_ (.A(_03068_),
    .B(_03069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03070_));
 sky130_fd_sc_hd__and2_2 _12136_ (.A(_02831_),
    .B(_02843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03071_));
 sky130_fd_sc_hd__a32o_2 _12137_ (.A1(_02832_),
    .A2(_02839_),
    .A3(_02840_),
    .B1(_02831_),
    .B2(_02843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03072_));
 sky130_fd_sc_hd__o211a_2 _12138_ (.A1(_02831_),
    .A2(_02844_),
    .B1(_03070_),
    .C1(_02843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03073_));
 sky130_fd_sc_hd__o2bb2ai_2 _12139_ (.A1_N(_03068_),
    .A2_N(_03069_),
    .B1(_03071_),
    .B2(_02844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03074_));
 sky130_fd_sc_hd__nor2_2 _12140_ (.A(_03070_),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03075_));
 sky130_fd_sc_hd__nand3b_2 _12141_ (.A_N(_03072_),
    .B(_03069_),
    .C(_03068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03076_));
 sky130_fd_sc_hd__a21o_2 _12142_ (.A1(_03068_),
    .A2(_03069_),
    .B1(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03077_));
 sky130_fd_sc_hd__nand2_2 _12143_ (.A(_03069_),
    .B(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03078_));
 sky130_fd_sc_hd__o2111ai_2 _12144_ (.A1(_02831_),
    .A2(_02844_),
    .B1(_03068_),
    .C1(_03069_),
    .D1(_02843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_2 _12145_ (.A(_03077_),
    .B(_03079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2_2 _12146_ (.A(_03074_),
    .B(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03081_));
 sky130_fd_sc_hd__nand4_2 _12147_ (.A(_03035_),
    .B(_03037_),
    .C(_03074_),
    .D(_03076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03082_));
 sky130_fd_sc_hd__o2bb2ai_2 _12148_ (.A1_N(_03035_),
    .A2_N(_03037_),
    .B1(_03073_),
    .B2(_03075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03083_));
 sky130_fd_sc_hd__a21oi_2 _12149_ (.A1(_03035_),
    .A2(_03037_),
    .B1(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03084_));
 sky130_fd_sc_hd__nand3_2 _12150_ (.A(_03035_),
    .B(_03037_),
    .C(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_2 _12151_ (.A(_02925_),
    .B(_02858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03086_));
 sky130_fd_sc_hd__o2bb2ai_2 _12152_ (.A1_N(_02858_),
    .A2_N(_02925_),
    .B1(_02927_),
    .B2(_02922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03087_));
 sky130_fd_sc_hd__nand3_2 _12153_ (.A(_03087_),
    .B(_03083_),
    .C(_03082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03088_));
 sky130_fd_sc_hd__nand3_2 _12154_ (.A(_02928_),
    .B(_03085_),
    .C(_03086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03089_));
 sky130_fd_sc_hd__o21ai_2 _12155_ (.A1(_03084_),
    .A2(_03089_),
    .B1(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03090_));
 sky130_fd_sc_hd__a21bo_2 _12156_ (.A1(_02829_),
    .A2(_02827_),
    .B1_N(_02828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03091_));
 sky130_fd_sc_hd__a31o_2 _12157_ (.A1(_02825_),
    .A2(_02847_),
    .A3(_02848_),
    .B1(_02854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03092_));
 sky130_fd_sc_hd__and3_2 _12158_ (.A(_02852_),
    .B(_03091_),
    .C(_03092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03093_));
 sky130_fd_sc_hd__nand3_2 _12159_ (.A(_02852_),
    .B(_03091_),
    .C(_03092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03094_));
 sky130_fd_sc_hd__nand3b_2 _12160_ (.A_N(_03091_),
    .B(_02856_),
    .C(_02851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03095_));
 sky130_fd_sc_hd__a22oi_2 _12161_ (.A1(\a_h[1] ),
    .A2(\b_h[15] ),
    .B1(_03094_),
    .B2(_03095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03096_));
 sky130_fd_sc_hd__and4_2 _12162_ (.A(_03094_),
    .B(_03095_),
    .C(\a_h[1] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03097_));
 sky130_fd_sc_hd__nor2_2 _12163_ (.A(_03096_),
    .B(_03097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03098_));
 sky130_fd_sc_hd__nand2_2 _12164_ (.A(_03090_),
    .B(_03098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03099_));
 sky130_fd_sc_hd__o221ai_2 _12165_ (.A1(_03096_),
    .A2(_03097_),
    .B1(_03084_),
    .B2(_03089_),
    .C1(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03100_));
 sky130_fd_sc_hd__o211a_2 _12166_ (.A1(_03084_),
    .A2(_03089_),
    .B1(_03098_),
    .C1(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03101_));
 sky130_fd_sc_hd__o211ai_2 _12167_ (.A1(_03084_),
    .A2(_03089_),
    .B1(_03098_),
    .C1(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03102_));
 sky130_fd_sc_hd__o21ai_2 _12168_ (.A1(_03096_),
    .A2(_03097_),
    .B1(_03090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03103_));
 sky130_fd_sc_hd__nand3_2 _12169_ (.A(_02967_),
    .B(_03099_),
    .C(_03100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_2 _12170_ (.A(_02968_),
    .B(_03103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03105_));
 sky130_fd_sc_hd__nand3_2 _12171_ (.A(_02968_),
    .B(_03102_),
    .C(_03103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03106_));
 sky130_fd_sc_hd__nor3_2 _12172_ (.A(_09177_),
    .B(_09679_),
    .C(_02941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03107_));
 sky130_fd_sc_hd__a31o_2 _12173_ (.A1(_02789_),
    .A2(_02938_),
    .A3(_02939_),
    .B1(_03107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03108_));
 sky130_fd_sc_hd__inv_2 _12174_ (.A(_03108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03109_));
 sky130_fd_sc_hd__o2bb2ai_2 _12175_ (.A1_N(_03104_),
    .A2_N(_03106_),
    .B1(_03107_),
    .B2(_02940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03110_));
 sky130_fd_sc_hd__nand3_2 _12176_ (.A(_03104_),
    .B(_03106_),
    .C(_03109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_2 _12177_ (.A(_03110_),
    .B(_03111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03112_));
 sky130_fd_sc_hd__a2bb2o_2 _12178_ (.A1_N(_02949_),
    .A2_N(_02952_),
    .B1(_02695_),
    .B2(_02955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03113_));
 sky130_fd_sc_hd__nand4_2 _12179_ (.A(_02954_),
    .B(_02957_),
    .C(_03110_),
    .D(_03111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03114_));
 sky130_fd_sc_hd__nand2_2 _12180_ (.A(_03112_),
    .B(_03113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03115_));
 sky130_fd_sc_hd__and2_2 _12181_ (.A(_03114_),
    .B(_03115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03116_));
 sky130_fd_sc_hd__o21ai_2 _12182_ (.A1(_02813_),
    .A2(_02962_),
    .B1(_02959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03117_));
 sky130_fd_sc_hd__o21a_2 _12183_ (.A1(_02688_),
    .A2(_02811_),
    .B1(_02959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03118_));
 sky130_fd_sc_hd__nand3_2 _12184_ (.A(_02817_),
    .B(_02818_),
    .C(_03118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03119_));
 sky130_fd_sc_hd__a22oi_2 _12185_ (.A1(_02815_),
    .A2(_02816_),
    .B1(_02963_),
    .B2(_02812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03120_));
 sky130_fd_sc_hd__nand3_2 _12186_ (.A(_03120_),
    .B(_02959_),
    .C(_02818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03121_));
 sky130_fd_sc_hd__a21oi_2 _12187_ (.A1(_03119_),
    .A2(_03117_),
    .B1(_03116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03122_));
 sky130_fd_sc_hd__and3_2 _12188_ (.A(_03119_),
    .B(_03117_),
    .C(_03116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03123_));
 sky130_fd_sc_hd__a311oi_2 _12189_ (.A1(_03116_),
    .A2(_03119_),
    .A3(_03117_),
    .B1(rst),
    .C1(_03122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00290_));
 sky130_fd_sc_hd__a22oi_2 _12190_ (.A1(_03036_),
    .A2(_03032_),
    .B1(_03035_),
    .B2(_03081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03124_));
 sky130_fd_sc_hd__a21oi_2 _12191_ (.A1(_03037_),
    .A2(_03080_),
    .B1(_03034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03125_));
 sky130_fd_sc_hd__a21o_2 _12192_ (.A1(_03006_),
    .A2(_03009_),
    .B1(_03010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03126_));
 sky130_fd_sc_hd__a21oi_2 _12193_ (.A1(_03006_),
    .A2(_03009_),
    .B1(_03010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03127_));
 sky130_fd_sc_hd__nand2_2 _12194_ (.A(\a_h[11] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03128_));
 sky130_fd_sc_hd__a22oi_2 _12195_ (.A1(\a_h[11] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_2 _12196_ (.A(_02978_),
    .B(_03128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_2 _12197_ (.A(\a_h[11] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03131_));
 sky130_fd_sc_hd__nand4_2 _12198_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03132_));
 sky130_fd_sc_hd__nand2_2 _12199_ (.A(\a_h[9] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03133_));
 sky130_fd_sc_hd__o2bb2ai_2 _12200_ (.A1_N(_03130_),
    .A2_N(_03132_),
    .B1(_09471_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03134_));
 sky130_fd_sc_hd__o2111ai_2 _12201_ (.A1(_02976_),
    .A2(_03131_),
    .B1(\a_h[9] ),
    .C1(\b_h[8] ),
    .D1(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03135_));
 sky130_fd_sc_hd__a21o_2 _12202_ (.A1(_03130_),
    .A2(_03132_),
    .B1(_03133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03136_));
 sky130_fd_sc_hd__o221ai_2 _12203_ (.A1(_09471_),
    .A2(_09613_),
    .B1(_02976_),
    .B2(_03131_),
    .C1(_03130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03137_));
 sky130_fd_sc_hd__nand3_2 _12204_ (.A(_03136_),
    .B(_03137_),
    .C(_03126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03138_));
 sky130_fd_sc_hd__nand3_2 _12205_ (.A(_03127_),
    .B(_03134_),
    .C(_03135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03139_));
 sky130_fd_sc_hd__a22oi_2 _12206_ (.A1(_02864_),
    .A2(_02976_),
    .B1(_02979_),
    .B2(_02975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03140_));
 sky130_fd_sc_hd__inv_2 _12207_ (.A(_03140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03141_));
 sky130_fd_sc_hd__a21o_2 _12208_ (.A1(_03138_),
    .A2(_03139_),
    .B1(_03140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03142_));
 sky130_fd_sc_hd__nand3_2 _12209_ (.A(_03138_),
    .B(_03139_),
    .C(_03140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03143_));
 sky130_fd_sc_hd__nand3_2 _12210_ (.A(_03138_),
    .B(_03139_),
    .C(_03141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03144_));
 sky130_fd_sc_hd__a21o_2 _12211_ (.A1(_03138_),
    .A2(_03139_),
    .B1(_03141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03145_));
 sky130_fd_sc_hd__nand2_2 _12212_ (.A(_03144_),
    .B(_03145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03146_));
 sky130_fd_sc_hd__and3_2 _12213_ (.A(_02738_),
    .B(\b_h[2] ),
    .C(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03147_));
 sky130_fd_sc_hd__nand2_2 _12214_ (.A(\a_h[12] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2_2 _12215_ (.A(\a_h[14] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_2 _12216_ (.A(_03007_),
    .B(_03149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03150_));
 sky130_fd_sc_hd__nand2_2 _12217_ (.A(\a_h[14] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03151_));
 sky130_fd_sc_hd__nand4_2 _12218_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03152_));
 sky130_fd_sc_hd__o221ai_2 _12219_ (.A1(_09504_),
    .A2(_09602_),
    .B1(_03008_),
    .B2(_03151_),
    .C1(_03150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03153_));
 sky130_fd_sc_hd__a21o_2 _12220_ (.A1(_03150_),
    .A2(_03152_),
    .B1(_03148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03154_));
 sky130_fd_sc_hd__o2111ai_2 _12221_ (.A1(_03008_),
    .A2(_03151_),
    .B1(\a_h[12] ),
    .C1(\b_h[5] ),
    .D1(_03150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03155_));
 sky130_fd_sc_hd__a21bo_2 _12222_ (.A1(_03150_),
    .A2(_03152_),
    .B1_N(_03148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03156_));
 sky130_fd_sc_hd__nand3_2 _12223_ (.A(_03156_),
    .B(_03147_),
    .C(_03155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03157_));
 sky130_fd_sc_hd__inv_2 _12224_ (.A(_03157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03158_));
 sky130_fd_sc_hd__nand3b_2 _12225_ (.A_N(_03147_),
    .B(_03153_),
    .C(_03154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_2 _12226_ (.A(_03157_),
    .B(_03159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03160_));
 sky130_fd_sc_hd__o21a_2 _12227_ (.A1(_03004_),
    .A2(_03022_),
    .B1(_03160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03161_));
 sky130_fd_sc_hd__o21ai_2 _12228_ (.A1(_03004_),
    .A2(_03022_),
    .B1(_03160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03162_));
 sky130_fd_sc_hd__nand4_2 _12229_ (.A(_03003_),
    .B(_03023_),
    .C(_03157_),
    .D(_03159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_2 _12230_ (.A(_03162_),
    .B(_03163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03164_));
 sky130_fd_sc_hd__nand4_2 _12231_ (.A(_03144_),
    .B(_03145_),
    .C(_03162_),
    .D(_03163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_2 _12232_ (.A(_03164_),
    .B(_03146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03166_));
 sky130_fd_sc_hd__a22o_2 _12233_ (.A1(_03142_),
    .A2(_03143_),
    .B1(_03162_),
    .B2(_03163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03167_));
 sky130_fd_sc_hd__nand4_2 _12234_ (.A(_03142_),
    .B(_03143_),
    .C(_03162_),
    .D(_03163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03168_));
 sky130_fd_sc_hd__nand4_2 _12235_ (.A(_03026_),
    .B(_03028_),
    .C(_03165_),
    .D(_03166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03169_));
 sky130_fd_sc_hd__a22oi_2 _12236_ (.A1(_03026_),
    .A2(_03028_),
    .B1(_03165_),
    .B2(_03166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03170_));
 sky130_fd_sc_hd__nand3_2 _12237_ (.A(_03033_),
    .B(_03167_),
    .C(_03168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_2 _12238_ (.A(_03169_),
    .B(_03171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03172_));
 sky130_fd_sc_hd__a31oi_2 _12239_ (.A1(_02973_),
    .A2(_02981_),
    .A3(_02982_),
    .B1(_02990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03173_));
 sky130_fd_sc_hd__a21o_2 _12240_ (.A1(_02986_),
    .A2(_02990_),
    .B1(_02987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03174_));
 sky130_fd_sc_hd__nand2_2 _12241_ (.A(\a_h[5] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03175_));
 sky130_fd_sc_hd__a22o_2 _12242_ (.A1(\a_h[5] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03176_));
 sky130_fd_sc_hd__a21o_2 _12243_ (.A1(\a_h[5] ),
    .A2(\b_h[12] ),
    .B1(_03043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03177_));
 sky130_fd_sc_hd__o2111a_2 _12244_ (.A1(_03041_),
    .A2(_03175_),
    .B1(\a_h[3] ),
    .C1(\b_h[14] ),
    .D1(_03176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03178_));
 sky130_fd_sc_hd__a32oi_2 _12245_ (.A1(_03043_),
    .A2(\b_h[12] ),
    .A3(\a_h[5] ),
    .B1(\a_h[3] ),
    .B2(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03179_));
 sky130_fd_sc_hd__a21oi_2 _12246_ (.A1(_03177_),
    .A2(_03179_),
    .B1(_03178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03180_));
 sky130_fd_sc_hd__a21o_2 _12247_ (.A1(_03177_),
    .A2(_03179_),
    .B1(_03178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03181_));
 sky130_fd_sc_hd__o21ai_2 _12248_ (.A1(_03050_),
    .A2(_03052_),
    .B1(_03055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03182_));
 sky130_fd_sc_hd__o22a_2 _12249_ (.A1(_02833_),
    .A2(_03054_),
    .B1(_03050_),
    .B2(_03052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03183_));
 sky130_fd_sc_hd__nand2_2 _12250_ (.A(\a_h[8] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03184_));
 sky130_fd_sc_hd__a22oi_2 _12251_ (.A1(\a_h[8] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_2 _12252_ (.A(_03054_),
    .B(_03184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03186_));
 sky130_fd_sc_hd__nand4_2 _12253_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_2 _12254_ (.A(\a_h[6] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03188_));
 sky130_fd_sc_hd__a21o_2 _12255_ (.A1(_03186_),
    .A2(_03187_),
    .B1(_03188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03189_));
 sky130_fd_sc_hd__o211ai_2 _12256_ (.A1(_09439_),
    .A2(_09646_),
    .B1(_03186_),
    .C1(_03187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03190_));
 sky130_fd_sc_hd__nand4_2 _12257_ (.A(_03186_),
    .B(_03187_),
    .C(\a_h[6] ),
    .D(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03191_));
 sky130_fd_sc_hd__a22o_2 _12258_ (.A1(\a_h[6] ),
    .A2(\b_h[11] ),
    .B1(_03186_),
    .B2(_03187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03192_));
 sky130_fd_sc_hd__and3_2 _12259_ (.A(_03192_),
    .B(_03182_),
    .C(_03191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03193_));
 sky130_fd_sc_hd__nand3_2 _12260_ (.A(_03192_),
    .B(_03182_),
    .C(_03191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03194_));
 sky130_fd_sc_hd__nand3_2 _12261_ (.A(_03183_),
    .B(_03189_),
    .C(_03190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03195_));
 sky130_fd_sc_hd__nand2_2 _12262_ (.A(_03194_),
    .B(_03195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_2 _12263_ (.A(_03180_),
    .B(_03195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03197_));
 sky130_fd_sc_hd__a21o_2 _12264_ (.A1(_03194_),
    .A2(_03195_),
    .B1(_03180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03198_));
 sky130_fd_sc_hd__nand3_2 _12265_ (.A(_03181_),
    .B(_03194_),
    .C(_03195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03199_));
 sky130_fd_sc_hd__nand2_2 _12266_ (.A(_03196_),
    .B(_03180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03200_));
 sky130_fd_sc_hd__o211ai_2 _12267_ (.A1(_03193_),
    .A2(_03197_),
    .B1(_03174_),
    .C1(_03198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03201_));
 sky130_fd_sc_hd__o211ai_2 _12268_ (.A1(_02985_),
    .A2(_03173_),
    .B1(_03199_),
    .C1(_03200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03202_));
 sky130_fd_sc_hd__o31a_2 _12269_ (.A1(_03045_),
    .A2(_03046_),
    .A3(_03060_),
    .B1(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03203_));
 sky130_fd_sc_hd__o31ai_2 _12270_ (.A1(_03045_),
    .A2(_03046_),
    .A3(_03060_),
    .B1(_03062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03204_));
 sky130_fd_sc_hd__and3_2 _12271_ (.A(_03201_),
    .B(_03202_),
    .C(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03205_));
 sky130_fd_sc_hd__nand3_2 _12272_ (.A(_03201_),
    .B(_03202_),
    .C(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03206_));
 sky130_fd_sc_hd__a21oi_2 _12273_ (.A1(_03201_),
    .A2(_03202_),
    .B1(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03207_));
 sky130_fd_sc_hd__a21o_2 _12274_ (.A1(_03201_),
    .A2(_03202_),
    .B1(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03208_));
 sky130_fd_sc_hd__a22o_2 _12275_ (.A1(_03061_),
    .A2(_03066_),
    .B1(_03201_),
    .B2(_03202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03209_));
 sky130_fd_sc_hd__nand2_2 _12276_ (.A(_03202_),
    .B(_03204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03210_));
 sky130_fd_sc_hd__nand4_2 _12277_ (.A(_03061_),
    .B(_03066_),
    .C(_03201_),
    .D(_03202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_2 _12278_ (.A(_03209_),
    .B(_03211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_2 _12279_ (.A(_03206_),
    .B(_03208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03213_));
 sky130_fd_sc_hd__nand2_2 _12280_ (.A(_03172_),
    .B(_03212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03214_));
 sky130_fd_sc_hd__nand4_2 _12281_ (.A(_03169_),
    .B(_03171_),
    .C(_03209_),
    .D(_03211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03215_));
 sky130_fd_sc_hd__nand4_2 _12282_ (.A(_03169_),
    .B(_03171_),
    .C(_03206_),
    .D(_03208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03216_));
 sky130_fd_sc_hd__o2bb2ai_2 _12283_ (.A1_N(_03169_),
    .A2_N(_03171_),
    .B1(_03205_),
    .B2(_03207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03217_));
 sky130_fd_sc_hd__nand3_2 _12284_ (.A(_03125_),
    .B(_03214_),
    .C(_03215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03218_));
 sky130_fd_sc_hd__nand3_2 _12285_ (.A(_03124_),
    .B(_03216_),
    .C(_03217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_2 _12286_ (.A(_03218_),
    .B(_03219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03220_));
 sky130_fd_sc_hd__a31oi_2 _12287_ (.A1(\a_h[3] ),
    .A2(\a_h[4] ),
    .A3(_02588_),
    .B1(_03045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03221_));
 sky130_fd_sc_hd__a32oi_2 _12288_ (.A1(_03038_),
    .A2(_03064_),
    .A3(_03065_),
    .B1(_03069_),
    .B2(_03072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03222_));
 sky130_fd_sc_hd__a21oi_2 _12289_ (.A1(_03068_),
    .A2(_03078_),
    .B1(_03221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03223_));
 sky130_fd_sc_hd__and3_2 _12290_ (.A(_03068_),
    .B(_03078_),
    .C(_03221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03224_));
 sky130_fd_sc_hd__nand2_2 _12291_ (.A(_03221_),
    .B(_03222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03225_));
 sky130_fd_sc_hd__nor2_2 _12292_ (.A(_09395_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03226_));
 sky130_fd_sc_hd__o22a_2 _12293_ (.A1(_09395_),
    .A2(_09679_),
    .B1(_03221_),
    .B2(_03222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03227_));
 sky130_fd_sc_hd__o22ai_2 _12294_ (.A1(_09395_),
    .A2(_09679_),
    .B1(_03221_),
    .B2(_03222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03228_));
 sky130_fd_sc_hd__o21ai_2 _12295_ (.A1(_03223_),
    .A2(_03224_),
    .B1(_03226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03229_));
 sky130_fd_sc_hd__o21a_2 _12296_ (.A1(_03224_),
    .A2(_03228_),
    .B1(_03229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03230_));
 sky130_fd_sc_hd__o21ai_2 _12297_ (.A1(_03224_),
    .A2(_03228_),
    .B1(_03229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03231_));
 sky130_fd_sc_hd__o2111ai_2 _12298_ (.A1(_03224_),
    .A2(_03228_),
    .B1(_03229_),
    .C1(_03219_),
    .D1(_03218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03232_));
 sky130_fd_sc_hd__a21o_2 _12299_ (.A1(_03218_),
    .A2(_03219_),
    .B1(_03230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03233_));
 sky130_fd_sc_hd__nand3_2 _12300_ (.A(_03218_),
    .B(_03219_),
    .C(_03231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_2 _12301_ (.A(_03220_),
    .B(_03230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03235_));
 sky130_fd_sc_hd__o2bb2ai_2 _12302_ (.A1_N(_03098_),
    .A2_N(_03088_),
    .B1(_03084_),
    .B2(_03089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03236_));
 sky130_fd_sc_hd__a2bb2oi_2 _12303_ (.A1_N(_03084_),
    .A2_N(_03089_),
    .B1(_03098_),
    .B2(_03088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03237_));
 sky130_fd_sc_hd__nand3_2 _12304_ (.A(_03232_),
    .B(_03233_),
    .C(_03237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03238_));
 sky130_fd_sc_hd__nand3_2 _12305_ (.A(_03236_),
    .B(_03235_),
    .C(_03234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03239_));
 sky130_fd_sc_hd__a31o_2 _12306_ (.A1(\a_h[1] ),
    .A2(_03095_),
    .A3(\b_h[15] ),
    .B1(_03093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03240_));
 sky130_fd_sc_hd__a21oi_2 _12307_ (.A1(_03238_),
    .A2(_03239_),
    .B1(_03240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03241_));
 sky130_fd_sc_hd__a21o_2 _12308_ (.A1(_03238_),
    .A2(_03239_),
    .B1(_03240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03242_));
 sky130_fd_sc_hd__nand2_2 _12309_ (.A(_03238_),
    .B(_03240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03243_));
 sky130_fd_sc_hd__and3_2 _12310_ (.A(_03238_),
    .B(_03239_),
    .C(_03240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03244_));
 sky130_fd_sc_hd__o2bb2ai_2 _12311_ (.A1_N(_03108_),
    .A2_N(_03104_),
    .B1(_03101_),
    .B2(_03105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03245_));
 sky130_fd_sc_hd__a32o_2 _12312_ (.A1(_02967_),
    .A2(_03099_),
    .A3(_03100_),
    .B1(_03106_),
    .B2(_03109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03246_));
 sky130_fd_sc_hd__o21ai_2 _12313_ (.A1(_03241_),
    .A2(_03244_),
    .B1(_03246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_2 _12314_ (.A(_03242_),
    .B(_03245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03248_));
 sky130_fd_sc_hd__o21ai_2 _12315_ (.A1(_03244_),
    .A2(_03248_),
    .B1(_03247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03249_));
 sky130_fd_sc_hd__a21oi_2 _12316_ (.A1(_03112_),
    .A2(_03113_),
    .B1(_03123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03250_));
 sky130_fd_sc_hd__a21oi_2 _12317_ (.A1(_03250_),
    .A2(_03249_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03251_));
 sky130_fd_sc_hd__o21a_2 _12318_ (.A1(_03249_),
    .A2(_03250_),
    .B1(_03251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00291_));
 sky130_fd_sc_hd__a32oi_2 _12319_ (.A1(_03125_),
    .A2(_03214_),
    .A3(_03215_),
    .B1(_03219_),
    .B2(_03231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03252_));
 sky130_fd_sc_hd__o32a_2 _12320_ (.A1(_09471_),
    .A2(_09613_),
    .A3(_03129_),
    .B1(_03131_),
    .B2(_02976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03253_));
 sky130_fd_sc_hd__a21oi_2 _12321_ (.A1(_03132_),
    .A2(_03133_),
    .B1(_03129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03254_));
 sky130_fd_sc_hd__a22oi_2 _12322_ (.A1(_03007_),
    .A2(_03149_),
    .B1(_03152_),
    .B2(_03148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03255_));
 sky130_fd_sc_hd__a22o_2 _12323_ (.A1(_03007_),
    .A2(_03149_),
    .B1(_03152_),
    .B2(_03148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03256_));
 sky130_fd_sc_hd__nand2_2 _12324_ (.A(\a_h[10] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03257_));
 sky130_fd_sc_hd__nand2_2 _12325_ (.A(\a_h[12] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03258_));
 sky130_fd_sc_hd__a22oi_2 _12326_ (.A1(\a_h[12] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_2 _12327_ (.A(_03131_),
    .B(_03258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_2 _12328_ (.A(\a_h[12] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03261_));
 sky130_fd_sc_hd__and4_2 _12329_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03262_));
 sky130_fd_sc_hd__nand4_2 _12330_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03263_));
 sky130_fd_sc_hd__a22o_2 _12331_ (.A1(\a_h[10] ),
    .A2(\b_h[8] ),
    .B1(_03260_),
    .B2(_03263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03264_));
 sky130_fd_sc_hd__o2111ai_2 _12332_ (.A1(_03128_),
    .A2(_03261_),
    .B1(\a_h[10] ),
    .C1(\b_h[8] ),
    .D1(_03260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03265_));
 sky130_fd_sc_hd__o221ai_2 _12333_ (.A1(_09482_),
    .A2(_09613_),
    .B1(_03128_),
    .B2(_03261_),
    .C1(_03260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03266_));
 sky130_fd_sc_hd__a21o_2 _12334_ (.A1(_03260_),
    .A2(_03263_),
    .B1(_03257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03267_));
 sky130_fd_sc_hd__nand3_2 _12335_ (.A(_03256_),
    .B(_03266_),
    .C(_03267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03268_));
 sky130_fd_sc_hd__nand3_2 _12336_ (.A(_03264_),
    .B(_03265_),
    .C(_03255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03269_));
 sky130_fd_sc_hd__a32oi_2 _12337_ (.A1(_03256_),
    .A2(_03266_),
    .A3(_03267_),
    .B1(_03269_),
    .B2(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03270_));
 sky130_fd_sc_hd__a32o_2 _12338_ (.A1(_03256_),
    .A2(_03266_),
    .A3(_03267_),
    .B1(_03269_),
    .B2(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03271_));
 sky130_fd_sc_hd__a21oi_2 _12339_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_2 _12340_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03273_));
 sky130_fd_sc_hd__and3_2 _12341_ (.A(_03268_),
    .B(_03269_),
    .C(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03274_));
 sky130_fd_sc_hd__nand3_2 _12342_ (.A(_03268_),
    .B(_03269_),
    .C(_03253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03275_));
 sky130_fd_sc_hd__a21o_2 _12343_ (.A1(_03268_),
    .A2(_03269_),
    .B1(_03254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03276_));
 sky130_fd_sc_hd__nand3_2 _12344_ (.A(_03254_),
    .B(_03268_),
    .C(_03269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_2 _12345_ (.A(\a_h[13] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_2 _12346_ (.A(\a_h[15] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03279_));
 sky130_fd_sc_hd__nand4_2 _12347_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[3] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03280_));
 sky130_fd_sc_hd__a22oi_2 _12348_ (.A1(\a_h[15] ),
    .A2(\b_h[3] ),
    .B1(\b_h[4] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_2 _12349_ (.A(_03151_),
    .B(_03279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03282_));
 sky130_fd_sc_hd__and3_2 _12350_ (.A(_03278_),
    .B(_03280_),
    .C(_03282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03283_));
 sky130_fd_sc_hd__a21oi_2 _12351_ (.A1(_03280_),
    .A2(_03282_),
    .B1(_03278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03284_));
 sky130_fd_sc_hd__nor2_2 _12352_ (.A(_03283_),
    .B(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03285_));
 sky130_fd_sc_hd__o21ai_2 _12353_ (.A1(_02899_),
    .A2(_02996_),
    .B1(_03285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03286_));
 sky130_fd_sc_hd__o211ai_2 _12354_ (.A1(_02899_),
    .A2(_02996_),
    .B1(_03157_),
    .C1(_03285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03287_));
 sky130_fd_sc_hd__o2bb2ai_2 _12355_ (.A1_N(_02998_),
    .A2_N(_03157_),
    .B1(_03283_),
    .B2(_03284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03288_));
 sky130_fd_sc_hd__nand2_2 _12356_ (.A(_03287_),
    .B(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03289_));
 sky130_fd_sc_hd__nand3_2 _12357_ (.A(_03273_),
    .B(_03275_),
    .C(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03290_));
 sky130_fd_sc_hd__nand4_2 _12358_ (.A(_03273_),
    .B(_03275_),
    .C(_03287_),
    .D(_03288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03291_));
 sky130_fd_sc_hd__o21ai_2 _12359_ (.A1(_03272_),
    .A2(_03274_),
    .B1(_03289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03292_));
 sky130_fd_sc_hd__nand3_2 _12360_ (.A(_03142_),
    .B(_03143_),
    .C(_03162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03293_));
 sky130_fd_sc_hd__a31oi_2 _12361_ (.A1(_03144_),
    .A2(_03145_),
    .A3(_03163_),
    .B1(_03161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03294_));
 sky130_fd_sc_hd__nand4_2 _12362_ (.A(_03163_),
    .B(_03291_),
    .C(_03292_),
    .D(_03293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03295_));
 sky130_fd_sc_hd__o2111ai_2 _12363_ (.A1(_03158_),
    .A2(_03286_),
    .B1(_03288_),
    .C1(_03276_),
    .D1(_03277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03296_));
 sky130_fd_sc_hd__nand3_2 _12364_ (.A(_03273_),
    .B(_03275_),
    .C(_03289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03297_));
 sky130_fd_sc_hd__nand3_2 _12365_ (.A(_03294_),
    .B(_03296_),
    .C(_03297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_2 _12366_ (.A(_03295_),
    .B(_03298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03299_));
 sky130_fd_sc_hd__nand2_2 _12367_ (.A(\a_h[6] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03300_));
 sky130_fd_sc_hd__and4_2 _12368_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03301_));
 sky130_fd_sc_hd__nand4_2 _12369_ (.A(\a_h[5] ),
    .B(\a_h[6] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2_2 _12370_ (.A(_03175_),
    .B(_03300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03303_));
 sky130_fd_sc_hd__and4_2 _12371_ (.A(_03303_),
    .B(\b_h[14] ),
    .C(\a_h[4] ),
    .D(_03302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03304_));
 sky130_fd_sc_hd__o2bb2a_2 _12372_ (.A1_N(_03302_),
    .A2_N(_03303_),
    .B1(_09417_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03305_));
 sky130_fd_sc_hd__nor2_2 _12373_ (.A(_03304_),
    .B(_03305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03306_));
 sky130_fd_sc_hd__a21o_2 _12374_ (.A1(_03187_),
    .A2(_03188_),
    .B1(_03185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03307_));
 sky130_fd_sc_hd__a21oi_2 _12375_ (.A1(_03187_),
    .A2(_03188_),
    .B1(_03185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_2 _12376_ (.A(\a_h[7] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03309_));
 sky130_fd_sc_hd__nand2_2 _12377_ (.A(\a_h[8] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03310_));
 sky130_fd_sc_hd__nand2_2 _12378_ (.A(\a_h[9] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03311_));
 sky130_fd_sc_hd__a22oi_2 _12379_ (.A1(\a_h[9] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03312_));
 sky130_fd_sc_hd__nand2_2 _12380_ (.A(_03310_),
    .B(_03311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_2 _12381_ (.A(\a_h[9] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03314_));
 sky130_fd_sc_hd__nand4_2 _12382_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03315_));
 sky130_fd_sc_hd__o2bb2ai_2 _12383_ (.A1_N(_03313_),
    .A2_N(_03315_),
    .B1(_09449_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03316_));
 sky130_fd_sc_hd__nand3_2 _12384_ (.A(_03315_),
    .B(\b_h[11] ),
    .C(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03317_));
 sky130_fd_sc_hd__o22a_2 _12385_ (.A1(_09449_),
    .A2(_09646_),
    .B1(_03310_),
    .B2(_03311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03318_));
 sky130_fd_sc_hd__o21ai_2 _12386_ (.A1(_03310_),
    .A2(_03311_),
    .B1(_03309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03319_));
 sky130_fd_sc_hd__a21o_2 _12387_ (.A1(_03313_),
    .A2(_03315_),
    .B1(_03309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03320_));
 sky130_fd_sc_hd__o211ai_2 _12388_ (.A1(_03312_),
    .A2(_03319_),
    .B1(_03307_),
    .C1(_03320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03321_));
 sky130_fd_sc_hd__o211a_2 _12389_ (.A1(_03317_),
    .A2(_03312_),
    .B1(_03308_),
    .C1(_03316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03322_));
 sky130_fd_sc_hd__o211ai_2 _12390_ (.A1(_03317_),
    .A2(_03312_),
    .B1(_03308_),
    .C1(_03316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_2 _12391_ (.A(_03321_),
    .B(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03324_));
 sky130_fd_sc_hd__o21ai_2 _12392_ (.A1(_03304_),
    .A2(_03305_),
    .B1(_03324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03325_));
 sky130_fd_sc_hd__nand3_2 _12393_ (.A(_03306_),
    .B(_03321_),
    .C(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03326_));
 sky130_fd_sc_hd__o211ai_2 _12394_ (.A1(_03304_),
    .A2(_03305_),
    .B1(_03321_),
    .C1(_03323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_2 _12395_ (.A(_03324_),
    .B(_03306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03328_));
 sky130_fd_sc_hd__a32oi_2 _12396_ (.A1(_03126_),
    .A2(_03136_),
    .A3(_03137_),
    .B1(_03139_),
    .B2(_03141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03329_));
 sky130_fd_sc_hd__a21boi_2 _12397_ (.A1(_03138_),
    .A2(_03140_),
    .B1_N(_03139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03330_));
 sky130_fd_sc_hd__nand3_2 _12398_ (.A(_03327_),
    .B(_03328_),
    .C(_03330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03331_));
 sky130_fd_sc_hd__nand3_2 _12399_ (.A(_03325_),
    .B(_03326_),
    .C(_03329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_2 _12400_ (.A(_03194_),
    .B(_03197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03333_));
 sky130_fd_sc_hd__a22o_2 _12401_ (.A1(_03194_),
    .A2(_03197_),
    .B1(_03331_),
    .B2(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03334_));
 sky130_fd_sc_hd__nand4_2 _12402_ (.A(_03194_),
    .B(_03197_),
    .C(_03331_),
    .D(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03335_));
 sky130_fd_sc_hd__a21oi_2 _12403_ (.A1(_03331_),
    .A2(_03332_),
    .B1(_03333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03336_));
 sky130_fd_sc_hd__a21o_2 _12404_ (.A1(_03331_),
    .A2(_03332_),
    .B1(_03333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03337_));
 sky130_fd_sc_hd__nand2_2 _12405_ (.A(_03331_),
    .B(_03333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03338_));
 sky130_fd_sc_hd__nand3_2 _12406_ (.A(_03331_),
    .B(_03332_),
    .C(_03333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03339_));
 sky130_fd_sc_hd__inv_2 _12407_ (.A(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03340_));
 sky130_fd_sc_hd__nand4_2 _12408_ (.A(_03295_),
    .B(_03298_),
    .C(_03334_),
    .D(_03335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03341_));
 sky130_fd_sc_hd__nand3_2 _12409_ (.A(_03299_),
    .B(_03337_),
    .C(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03342_));
 sky130_fd_sc_hd__nand4_2 _12410_ (.A(_03295_),
    .B(_03298_),
    .C(_03337_),
    .D(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03343_));
 sky130_fd_sc_hd__o2bb2ai_2 _12411_ (.A1_N(_03295_),
    .A2_N(_03298_),
    .B1(_03336_),
    .B2(_03340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03344_));
 sky130_fd_sc_hd__a31oi_2 _12412_ (.A1(_03169_),
    .A2(_03209_),
    .A3(_03211_),
    .B1(_03170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03345_));
 sky130_fd_sc_hd__nand3_2 _12413_ (.A(_03345_),
    .B(_03342_),
    .C(_03341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03346_));
 sky130_fd_sc_hd__o2111ai_2 _12414_ (.A1(_03170_),
    .A2(_03213_),
    .B1(_03343_),
    .C1(_03344_),
    .D1(_03169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03347_));
 sky130_fd_sc_hd__a41o_2 _12415_ (.A1(\a_h[4] ),
    .A2(\a_h[5] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_03178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03348_));
 sky130_fd_sc_hd__nand2_2 _12416_ (.A(_03201_),
    .B(_03203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03349_));
 sky130_fd_sc_hd__nand3_2 _12417_ (.A(_03202_),
    .B(_03348_),
    .C(_03349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03350_));
 sky130_fd_sc_hd__nand3b_2 _12418_ (.A_N(_03348_),
    .B(_03210_),
    .C(_03201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03351_));
 sky130_fd_sc_hd__a22o_2 _12419_ (.A1(\a_h[3] ),
    .A2(\b_h[15] ),
    .B1(_03350_),
    .B2(_03351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03352_));
 sky130_fd_sc_hd__nand4_2 _12420_ (.A(_03350_),
    .B(_03351_),
    .C(\a_h[3] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_2 _12421_ (.A(_03352_),
    .B(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03354_));
 sky130_fd_sc_hd__a22o_2 _12422_ (.A1(_03346_),
    .A2(_03347_),
    .B1(_03352_),
    .B2(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03355_));
 sky130_fd_sc_hd__nand4_2 _12423_ (.A(_03346_),
    .B(_03347_),
    .C(_03352_),
    .D(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03356_));
 sky130_fd_sc_hd__nand3b_2 _12424_ (.A_N(_03252_),
    .B(_03355_),
    .C(_03356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03357_));
 sky130_fd_sc_hd__nand3_2 _12425_ (.A(_03346_),
    .B(_03347_),
    .C(_03354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03358_));
 sky130_fd_sc_hd__a21o_2 _12426_ (.A1(_03346_),
    .A2(_03347_),
    .B1(_03354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03359_));
 sky130_fd_sc_hd__nand3_2 _12427_ (.A(_03359_),
    .B(_03252_),
    .C(_03358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03360_));
 sky130_fd_sc_hd__a31o_2 _12428_ (.A1(_03225_),
    .A2(\b_h[15] ),
    .A3(\a_h[2] ),
    .B1(_03223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03361_));
 sky130_fd_sc_hd__a21o_2 _12429_ (.A1(_03357_),
    .A2(_03360_),
    .B1(_03361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03362_));
 sky130_fd_sc_hd__nand2_2 _12430_ (.A(_03360_),
    .B(_03361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03363_));
 sky130_fd_sc_hd__nand4_2 _12431_ (.A(_03225_),
    .B(_03228_),
    .C(_03357_),
    .D(_03360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03364_));
 sky130_fd_sc_hd__a21bo_2 _12432_ (.A1(_03357_),
    .A2(_03360_),
    .B1_N(_03361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03365_));
 sky130_fd_sc_hd__o211ai_2 _12433_ (.A1(_03224_),
    .A2(_03227_),
    .B1(_03357_),
    .C1(_03360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03366_));
 sky130_fd_sc_hd__nand2_2 _12434_ (.A(_03239_),
    .B(_03243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03367_));
 sky130_fd_sc_hd__a21boi_2 _12435_ (.A1(_03238_),
    .A2(_03240_),
    .B1_N(_03239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03368_));
 sky130_fd_sc_hd__nand3_2 _12436_ (.A(_03365_),
    .B(_03366_),
    .C(_03368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03369_));
 sky130_fd_sc_hd__nand3_2 _12437_ (.A(_03362_),
    .B(_03367_),
    .C(_03364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03370_));
 sky130_fd_sc_hd__and2_2 _12438_ (.A(_03369_),
    .B(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03371_));
 sky130_fd_sc_hd__nand2_2 _12439_ (.A(_03369_),
    .B(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03372_));
 sky130_fd_sc_hd__o2bb2ai_2 _12440_ (.A1_N(_03112_),
    .A2_N(_03113_),
    .B1(_03244_),
    .B2(_03248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03373_));
 sky130_fd_sc_hd__o21ai_2 _12441_ (.A1(_03373_),
    .A2(_03123_),
    .B1(_03247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03374_));
 sky130_fd_sc_hd__o21ai_2 _12442_ (.A1(_03372_),
    .A2(_03374_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03375_));
 sky130_fd_sc_hd__a21oi_2 _12443_ (.A1(_03372_),
    .A2(_03374_),
    .B1(_03375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_2 _12444_ (.A(_03350_),
    .B(_03353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03376_));
 sky130_fd_sc_hd__inv_2 _12445_ (.A(_03376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03377_));
 sky130_fd_sc_hd__nand3_2 _12446_ (.A(_03298_),
    .B(_03334_),
    .C(_03335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03378_));
 sky130_fd_sc_hd__nand3_2 _12447_ (.A(_03295_),
    .B(_03337_),
    .C(_03339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_2 _12448_ (.A(_03298_),
    .B(_03379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03380_));
 sky130_fd_sc_hd__nand2_2 _12449_ (.A(_03295_),
    .B(_03378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03381_));
 sky130_fd_sc_hd__a21oi_2 _12450_ (.A1(_03309_),
    .A2(_03315_),
    .B1(_03312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03382_));
 sky130_fd_sc_hd__and2_2 _12451_ (.A(\a_h[8] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03383_));
 sky130_fd_sc_hd__nand2_2 _12452_ (.A(\a_h[8] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_2 _12453_ (.A(\a_h[10] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03385_));
 sky130_fd_sc_hd__a22oi_2 _12454_ (.A1(\a_h[10] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03386_));
 sky130_fd_sc_hd__nand2_2 _12455_ (.A(_03314_),
    .B(_03385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03387_));
 sky130_fd_sc_hd__nand3_2 _12456_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03388_));
 sky130_fd_sc_hd__nand4_2 _12457_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03389_));
 sky130_fd_sc_hd__a21oi_2 _12458_ (.A1(_03387_),
    .A2(_03389_),
    .B1(_03383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03390_));
 sky130_fd_sc_hd__a21o_2 _12459_ (.A1(_03387_),
    .A2(_03389_),
    .B1(_03383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03391_));
 sky130_fd_sc_hd__o211a_2 _12460_ (.A1(_09624_),
    .A2(_03388_),
    .B1(_03383_),
    .C1(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03392_));
 sky130_fd_sc_hd__o2111ai_2 _12461_ (.A1(_09624_),
    .A2(_03388_),
    .B1(\b_h[11] ),
    .C1(\a_h[8] ),
    .D1(_03387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03393_));
 sky130_fd_sc_hd__o22ai_2 _12462_ (.A1(_03312_),
    .A2(_03318_),
    .B1(_03390_),
    .B2(_03392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03394_));
 sky130_fd_sc_hd__nand3_2 _12463_ (.A(_03382_),
    .B(_03391_),
    .C(_03393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_2 _12464_ (.A(_03394_),
    .B(_03395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03396_));
 sky130_fd_sc_hd__nand2_2 _12465_ (.A(\a_h[7] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_2 _12466_ (.A(\a_h[6] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_2 _12467_ (.A(\a_h[7] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03399_));
 sky130_fd_sc_hd__nand2_2 _12468_ (.A(_03398_),
    .B(_03399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03400_));
 sky130_fd_sc_hd__a21o_2 _12469_ (.A1(\a_h[7] ),
    .A2(\b_h[12] ),
    .B1(_03398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03401_));
 sky130_fd_sc_hd__o2111a_2 _12470_ (.A1(_03300_),
    .A2(_03397_),
    .B1(\a_h[5] ),
    .C1(\b_h[14] ),
    .D1(_03400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03402_));
 sky130_fd_sc_hd__a32oi_2 _12471_ (.A1(_03398_),
    .A2(\b_h[12] ),
    .A3(\a_h[7] ),
    .B1(\a_h[5] ),
    .B2(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03403_));
 sky130_fd_sc_hd__a21oi_2 _12472_ (.A1(_03401_),
    .A2(_03403_),
    .B1(_03402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03404_));
 sky130_fd_sc_hd__a21o_2 _12473_ (.A1(_03401_),
    .A2(_03403_),
    .B1(_03402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03405_));
 sky130_fd_sc_hd__a21o_2 _12474_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_03404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03406_));
 sky130_fd_sc_hd__nand2_2 _12475_ (.A(_03404_),
    .B(_03394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03407_));
 sky130_fd_sc_hd__nand3_2 _12476_ (.A(_03394_),
    .B(_03404_),
    .C(_03395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03408_));
 sky130_fd_sc_hd__nand2_2 _12477_ (.A(_03396_),
    .B(_03404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03409_));
 sky130_fd_sc_hd__nand3_2 _12478_ (.A(_03394_),
    .B(_03395_),
    .C(_03405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03410_));
 sky130_fd_sc_hd__nand3_2 _12479_ (.A(_03271_),
    .B(_03409_),
    .C(_03410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03411_));
 sky130_fd_sc_hd__nand3_2 _12480_ (.A(_03406_),
    .B(_03408_),
    .C(_03270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03412_));
 sky130_fd_sc_hd__o21ai_2 _12481_ (.A1(_03306_),
    .A2(_03322_),
    .B1(_03321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03413_));
 sky130_fd_sc_hd__o21a_2 _12482_ (.A1(_03306_),
    .A2(_03322_),
    .B1(_03321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03414_));
 sky130_fd_sc_hd__a21o_2 _12483_ (.A1(_03411_),
    .A2(_03412_),
    .B1(_03414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03415_));
 sky130_fd_sc_hd__nand2_2 _12484_ (.A(_03411_),
    .B(_03414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03416_));
 sky130_fd_sc_hd__o2111ai_2 _12485_ (.A1(_03306_),
    .A2(_03322_),
    .B1(_03411_),
    .C1(_03412_),
    .D1(_03321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_2 _12486_ (.A(_03415_),
    .B(_03417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03418_));
 sky130_fd_sc_hd__and2_2 _12487_ (.A(\a_h[15] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03419_));
 sky130_fd_sc_hd__nand2_2 _12488_ (.A(\a_h[15] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03420_));
 sky130_fd_sc_hd__and4_2 _12489_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03421_));
 sky130_fd_sc_hd__or2_2 _12490_ (.A(_03151_),
    .B(_03420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03422_));
 sky130_fd_sc_hd__a22oi_2 _12491_ (.A1(\a_h[15] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03423_));
 sky130_fd_sc_hd__a22o_2 _12492_ (.A1(\a_h[15] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03424_));
 sky130_fd_sc_hd__a31o_2 _12493_ (.A1(\a_h[14] ),
    .A2(\b_h[4] ),
    .A3(_03419_),
    .B1(_03423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03425_));
 sky130_fd_sc_hd__o21a_2 _12494_ (.A1(_03151_),
    .A2(_03279_),
    .B1(_03278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03426_));
 sky130_fd_sc_hd__o21ai_2 _12495_ (.A1(_03278_),
    .A2(_03281_),
    .B1(_03280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03427_));
 sky130_fd_sc_hd__and2_2 _12496_ (.A(\a_h[11] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03428_));
 sky130_fd_sc_hd__nand2_2 _12497_ (.A(\a_h[11] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03429_));
 sky130_fd_sc_hd__nand2_2 _12498_ (.A(\a_h[13] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03430_));
 sky130_fd_sc_hd__a22o_2 _12499_ (.A1(\a_h[13] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_2 _12500_ (.A(\a_h[13] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03432_));
 sky130_fd_sc_hd__nand4_2 _12501_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03433_));
 sky130_fd_sc_hd__o2bb2ai_2 _12502_ (.A1_N(_03261_),
    .A2_N(_03430_),
    .B1(_03432_),
    .B2(_03258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03434_));
 sky130_fd_sc_hd__o21ai_2 _12503_ (.A1(_09493_),
    .A2(_09613_),
    .B1(_03434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03435_));
 sky130_fd_sc_hd__o211ai_2 _12504_ (.A1(_03258_),
    .A2(_03432_),
    .B1(_03428_),
    .C1(_03431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03436_));
 sky130_fd_sc_hd__o221ai_2 _12505_ (.A1(_09493_),
    .A2(_09613_),
    .B1(_03258_),
    .B2(_03432_),
    .C1(_03431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03437_));
 sky130_fd_sc_hd__nand2_2 _12506_ (.A(_03434_),
    .B(_03428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03438_));
 sky130_fd_sc_hd__o211ai_2 _12507_ (.A1(_03281_),
    .A2(_03426_),
    .B1(_03437_),
    .C1(_03438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03439_));
 sky130_fd_sc_hd__nand3_2 _12508_ (.A(_03435_),
    .B(_03436_),
    .C(_03427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03440_));
 sky130_fd_sc_hd__and3_2 _12509_ (.A(_03260_),
    .B(\b_h[8] ),
    .C(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03441_));
 sky130_fd_sc_hd__o22a_2 _12510_ (.A1(_09482_),
    .A2(_09613_),
    .B1(_03128_),
    .B2(_03261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03442_));
 sky130_fd_sc_hd__a31o_2 _12511_ (.A1(\a_h[10] ),
    .A2(_03260_),
    .A3(\b_h[8] ),
    .B1(_03262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03443_));
 sky130_fd_sc_hd__a21oi_2 _12512_ (.A1(_03439_),
    .A2(_03440_),
    .B1(_03443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03444_));
 sky130_fd_sc_hd__o2bb2ai_2 _12513_ (.A1_N(_03439_),
    .A2_N(_03440_),
    .B1(_03442_),
    .B2(_03259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03445_));
 sky130_fd_sc_hd__o211a_2 _12514_ (.A1(_03262_),
    .A2(_03441_),
    .B1(_03440_),
    .C1(_03439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03446_));
 sky130_fd_sc_hd__o211ai_2 _12515_ (.A1(_03262_),
    .A2(_03441_),
    .B1(_03440_),
    .C1(_03439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_2 _12516_ (.A(_03445_),
    .B(_03447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03448_));
 sky130_fd_sc_hd__a22oi_2 _12517_ (.A1(_03422_),
    .A2(_03424_),
    .B1(_03445_),
    .B2(_03447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03449_));
 sky130_fd_sc_hd__o22ai_2 _12518_ (.A1(_03421_),
    .A2(_03423_),
    .B1(_03444_),
    .B2(_03446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03450_));
 sky130_fd_sc_hd__nor3_2 _12519_ (.A(_03425_),
    .B(_03444_),
    .C(_03446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03451_));
 sky130_fd_sc_hd__nand3b_2 _12520_ (.A_N(_03425_),
    .B(_03445_),
    .C(_03447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03452_));
 sky130_fd_sc_hd__o211ai_2 _12521_ (.A1(_03158_),
    .A2(_03286_),
    .B1(_03290_),
    .C1(_03450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03453_));
 sky130_fd_sc_hd__o211ai_2 _12522_ (.A1(_03286_),
    .A2(_03158_),
    .B1(_03452_),
    .C1(_03290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03454_));
 sky130_fd_sc_hd__and4_2 _12523_ (.A(_03287_),
    .B(_03290_),
    .C(_03450_),
    .D(_03452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03455_));
 sky130_fd_sc_hd__o2bb2ai_2 _12524_ (.A1_N(_03287_),
    .A2_N(_03290_),
    .B1(_03449_),
    .B2(_03451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03456_));
 sky130_fd_sc_hd__o21ai_2 _12525_ (.A1(_03451_),
    .A2(_03453_),
    .B1(_03456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_2 _12526_ (.A(_03418_),
    .B(_03457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03458_));
 sky130_fd_sc_hd__o2111ai_2 _12527_ (.A1(_03449_),
    .A2(_03454_),
    .B1(_03456_),
    .C1(_03417_),
    .D1(_03415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03459_));
 sky130_fd_sc_hd__o211ai_2 _12528_ (.A1(_03451_),
    .A2(_03453_),
    .B1(_03456_),
    .C1(_03418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03460_));
 sky130_fd_sc_hd__nand3_2 _12529_ (.A(_03415_),
    .B(_03417_),
    .C(_03457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03461_));
 sky130_fd_sc_hd__a22oi_2 _12530_ (.A1(_03295_),
    .A2(_03378_),
    .B1(_03458_),
    .B2(_03459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03462_));
 sky130_fd_sc_hd__nand3_2 _12531_ (.A(_03381_),
    .B(_03460_),
    .C(_03461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03463_));
 sky130_fd_sc_hd__nand3_2 _12532_ (.A(_03380_),
    .B(_03458_),
    .C(_03459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03464_));
 sky130_fd_sc_hd__nor2_2 _12533_ (.A(_09417_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03465_));
 sky130_fd_sc_hd__nand2_2 _12534_ (.A(\a_h[4] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03466_));
 sky130_fd_sc_hd__a31o_2 _12535_ (.A1(\a_h[4] ),
    .A2(_03303_),
    .A3(\b_h[14] ),
    .B1(_03301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03467_));
 sky130_fd_sc_hd__nand3_2 _12536_ (.A(_03194_),
    .B(_03197_),
    .C(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03468_));
 sky130_fd_sc_hd__o211ai_2 _12537_ (.A1(_03301_),
    .A2(_03304_),
    .B1(_03331_),
    .C1(_03468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03469_));
 sky130_fd_sc_hd__nand3b_2 _12538_ (.A_N(_03467_),
    .B(_03338_),
    .C(_03332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03470_));
 sky130_fd_sc_hd__a31oi_2 _12539_ (.A1(_03331_),
    .A2(_03467_),
    .A3(_03468_),
    .B1(_03466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03471_));
 sky130_fd_sc_hd__and3_2 _12540_ (.A(_03469_),
    .B(_03470_),
    .C(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03472_));
 sky130_fd_sc_hd__nand2_2 _12541_ (.A(_03471_),
    .B(_03470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03473_));
 sky130_fd_sc_hd__a21oi_2 _12542_ (.A1(_03469_),
    .A2(_03470_),
    .B1(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03474_));
 sky130_fd_sc_hd__a21o_2 _12543_ (.A1(_03469_),
    .A2(_03470_),
    .B1(_03465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03475_));
 sky130_fd_sc_hd__a21oi_2 _12544_ (.A1(_03470_),
    .A2(_03471_),
    .B1(_03474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_2 _12545_ (.A(_03473_),
    .B(_03475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03477_));
 sky130_fd_sc_hd__a21oi_2 _12546_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03478_));
 sky130_fd_sc_hd__o2bb2ai_2 _12547_ (.A1_N(_03463_),
    .A2_N(_03464_),
    .B1(_03472_),
    .B2(_03474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03479_));
 sky130_fd_sc_hd__nand3_2 _12548_ (.A(_03463_),
    .B(_03464_),
    .C(_03476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_2 _12549_ (.A(_03347_),
    .B(_03354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03481_));
 sky130_fd_sc_hd__a21boi_2 _12550_ (.A1(_03347_),
    .A2(_03354_),
    .B1_N(_03346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03482_));
 sky130_fd_sc_hd__a21oi_2 _12551_ (.A1(_03479_),
    .A2(_03480_),
    .B1(_03482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03483_));
 sky130_fd_sc_hd__a21o_2 _12552_ (.A1(_03479_),
    .A2(_03480_),
    .B1(_03482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03484_));
 sky130_fd_sc_hd__nand3_2 _12553_ (.A(_03346_),
    .B(_03480_),
    .C(_03481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03485_));
 sky130_fd_sc_hd__nor2_2 _12554_ (.A(_03478_),
    .B(_03485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03486_));
 sky130_fd_sc_hd__o21ai_2 _12555_ (.A1(_03478_),
    .A2(_03485_),
    .B1(_03484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03487_));
 sky130_fd_sc_hd__o21ai_2 _12556_ (.A1(_03483_),
    .A2(_03486_),
    .B1(_03377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03488_));
 sky130_fd_sc_hd__o211ai_2 _12557_ (.A1(_03485_),
    .A2(_03478_),
    .B1(_03376_),
    .C1(_03484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_2 _12558_ (.A(_03357_),
    .B(_03363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03490_));
 sky130_fd_sc_hd__a21oi_2 _12559_ (.A1(_03488_),
    .A2(_03489_),
    .B1(_03490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03491_));
 sky130_fd_sc_hd__a21o_2 _12560_ (.A1(_03488_),
    .A2(_03489_),
    .B1(_03490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03492_));
 sky130_fd_sc_hd__a22oi_2 _12561_ (.A1(_03357_),
    .A2(_03363_),
    .B1(_03377_),
    .B2(_03487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03493_));
 sky130_fd_sc_hd__nand3_2 _12562_ (.A(_03488_),
    .B(_03489_),
    .C(_03490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03494_));
 sky130_fd_sc_hd__a21oi_2 _12563_ (.A1(_03493_),
    .A2(_03489_),
    .B1(_03491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_2 _12564_ (.A(_03492_),
    .B(_03494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03496_));
 sky130_fd_sc_hd__o21ai_2 _12565_ (.A1(_03372_),
    .A2(_03374_),
    .B1(_03370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03497_));
 sky130_fd_sc_hd__a21oi_2 _12566_ (.A1(_03497_),
    .A2(_03495_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03498_));
 sky130_fd_sc_hd__o21a_2 _12567_ (.A1(_03495_),
    .A2(_03497_),
    .B1(_03498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00293_));
 sky130_fd_sc_hd__o22a_2 _12568_ (.A1(_03485_),
    .A2(_03478_),
    .B1(_03377_),
    .B2(_03483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03499_));
 sky130_fd_sc_hd__a21bo_2 _12569_ (.A1(_03465_),
    .A2(_03470_),
    .B1_N(_03469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03500_));
 sky130_fd_sc_hd__a21boi_2 _12570_ (.A1(_03463_),
    .A2(_03476_),
    .B1_N(_03464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03501_));
 sky130_fd_sc_hd__o21ai_2 _12571_ (.A1(_03477_),
    .A2(_03462_),
    .B1(_03464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03502_));
 sky130_fd_sc_hd__a31oi_2 _12572_ (.A1(_03415_),
    .A2(_03417_),
    .A3(_03456_),
    .B1(_03455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03503_));
 sky130_fd_sc_hd__a31o_2 _12573_ (.A1(_03415_),
    .A2(_03417_),
    .A3(_03456_),
    .B1(_03455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03504_));
 sky130_fd_sc_hd__nand2_2 _12574_ (.A(\a_h[14] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_2 _12575_ (.A(_03432_),
    .B(_03505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_2 _12576_ (.A(\a_h[14] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03507_));
 sky130_fd_sc_hd__nand4_2 _12577_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03508_));
 sky130_fd_sc_hd__o2bb2ai_2 _12578_ (.A1_N(_03432_),
    .A2_N(_03505_),
    .B1(_03507_),
    .B2(_03430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03509_));
 sky130_fd_sc_hd__nand3_2 _12579_ (.A(_03506_),
    .B(_03508_),
    .C(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03510_));
 sky130_fd_sc_hd__nand4_2 _12580_ (.A(_03506_),
    .B(_03508_),
    .C(\a_h[12] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03511_));
 sky130_fd_sc_hd__o21ai_2 _12581_ (.A1(_09504_),
    .A2(_09613_),
    .B1(_03509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03512_));
 sky130_fd_sc_hd__o21ai_2 _12582_ (.A1(_09504_),
    .A2(_03510_),
    .B1(_03512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03513_));
 sky130_fd_sc_hd__a2bb2oi_2 _12583_ (.A1_N(_03151_),
    .A2_N(_03420_),
    .B1(_03511_),
    .B2(_03512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03514_));
 sky130_fd_sc_hd__o2bb2ai_2 _12584_ (.A1_N(_03511_),
    .A2_N(_03512_),
    .B1(_03151_),
    .B2(_03420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03515_));
 sky130_fd_sc_hd__a22oi_2 _12585_ (.A1(_03261_),
    .A2(_03430_),
    .B1(_03433_),
    .B2(_03429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _12586_ (.A(_03516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03517_));
 sky130_fd_sc_hd__o211a_2 _12587_ (.A1(_09504_),
    .A2(_03510_),
    .B1(_03421_),
    .C1(_03512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03518_));
 sky130_fd_sc_hd__o211ai_2 _12588_ (.A1(_09504_),
    .A2(_03510_),
    .B1(_03421_),
    .C1(_03512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03519_));
 sky130_fd_sc_hd__a31oi_2 _12589_ (.A1(_03512_),
    .A2(_03421_),
    .A3(_03511_),
    .B1(_03516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_2 _12590_ (.A(_03515_),
    .B(_03519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03521_));
 sky130_fd_sc_hd__nand3_2 _12591_ (.A(_03515_),
    .B(_03516_),
    .C(_03519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03522_));
 sky130_fd_sc_hd__nor2_2 _12592_ (.A(_03514_),
    .B(_03520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03523_));
 sky130_fd_sc_hd__a21oi_2 _12593_ (.A1(_03515_),
    .A2(_03516_),
    .B1(_03518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03524_));
 sky130_fd_sc_hd__o21ai_2 _12594_ (.A1(_03514_),
    .A2(_03518_),
    .B1(_03517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03525_));
 sky130_fd_sc_hd__nand3_2 _12595_ (.A(_03515_),
    .B(_03517_),
    .C(_03519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03526_));
 sky130_fd_sc_hd__a21oi_2 _12596_ (.A1(_03521_),
    .A2(_03517_),
    .B1(_03420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03527_));
 sky130_fd_sc_hd__nand3_2 _12597_ (.A(_03525_),
    .B(_03419_),
    .C(_03522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03528_));
 sky130_fd_sc_hd__a21oi_2 _12598_ (.A1(_03513_),
    .A2(_03516_),
    .B1(_03419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_2 _12599_ (.A(_03526_),
    .B(_03529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03530_));
 sky130_fd_sc_hd__a22o_2 _12600_ (.A1(_03529_),
    .A2(_03526_),
    .B1(_03527_),
    .B2(_03522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03531_));
 sky130_fd_sc_hd__o2bb2ai_2 _12601_ (.A1_N(_03528_),
    .A2_N(_03530_),
    .B1(_03425_),
    .B2(_03448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03532_));
 sky130_fd_sc_hd__nand3_2 _12602_ (.A(_03451_),
    .B(_03528_),
    .C(_03530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_2 _12603_ (.A(_03532_),
    .B(_03533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03534_));
 sky130_fd_sc_hd__a21boi_2 _12604_ (.A1(_03439_),
    .A2(_03443_),
    .B1_N(_03440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_2 _12605_ (.A(\a_h[9] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_2 _12606_ (.A(\a_h[10] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03537_));
 sky130_fd_sc_hd__nand2_2 _12607_ (.A(\a_h[11] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03538_));
 sky130_fd_sc_hd__nand4_2 _12608_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03539_));
 sky130_fd_sc_hd__a22oi_2 _12609_ (.A1(\a_h[11] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03540_));
 sky130_fd_sc_hd__nand2_2 _12610_ (.A(_03537_),
    .B(_03538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03541_));
 sky130_fd_sc_hd__o2bb2ai_2 _12611_ (.A1_N(_03539_),
    .A2_N(_03541_),
    .B1(_09471_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03542_));
 sky130_fd_sc_hd__nand4_2 _12612_ (.A(_03541_),
    .B(\b_h[11] ),
    .C(\a_h[9] ),
    .D(_03539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03543_));
 sky130_fd_sc_hd__o211ai_2 _12613_ (.A1(_09471_),
    .A2(_09646_),
    .B1(_03539_),
    .C1(_03541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03544_));
 sky130_fd_sc_hd__a21o_2 _12614_ (.A1(_03539_),
    .A2(_03541_),
    .B1(_03536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03545_));
 sky130_fd_sc_hd__a21oi_2 _12615_ (.A1(_03384_),
    .A2(_03389_),
    .B1(_03386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03546_));
 sky130_fd_sc_hd__a21oi_2 _12616_ (.A1(_03542_),
    .A2(_03543_),
    .B1(_03546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03547_));
 sky130_fd_sc_hd__nand3b_2 _12617_ (.A_N(_03546_),
    .B(_03545_),
    .C(_03544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03548_));
 sky130_fd_sc_hd__nand3_2 _12618_ (.A(_03542_),
    .B(_03543_),
    .C(_03546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_2 _12619_ (.A(\a_h[8] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03550_));
 sky130_fd_sc_hd__nand4_2 _12620_ (.A(\a_h[7] ),
    .B(\a_h[8] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03551_));
 sky130_fd_sc_hd__nand2_2 _12621_ (.A(_03397_),
    .B(_03550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2_2 _12622_ (.A(\a_h[6] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03553_));
 sky130_fd_sc_hd__nand4_2 _12623_ (.A(_03552_),
    .B(\b_h[14] ),
    .C(\a_h[6] ),
    .D(_03551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03554_));
 sky130_fd_sc_hd__o211ai_2 _12624_ (.A1(_09439_),
    .A2(_09668_),
    .B1(_03551_),
    .C1(_03552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03555_));
 sky130_fd_sc_hd__a21o_2 _12625_ (.A1(_03551_),
    .A2(_03552_),
    .B1(_03553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03556_));
 sky130_fd_sc_hd__nand2_2 _12626_ (.A(_03555_),
    .B(_03556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03557_));
 sky130_fd_sc_hd__a21oi_2 _12627_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03558_));
 sky130_fd_sc_hd__a21o_2 _12628_ (.A1(_03548_),
    .A2(_03549_),
    .B1(_03557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03559_));
 sky130_fd_sc_hd__and3_2 _12629_ (.A(_03548_),
    .B(_03557_),
    .C(_03549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03560_));
 sky130_fd_sc_hd__nand3_2 _12630_ (.A(_03548_),
    .B(_03557_),
    .C(_03549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03561_));
 sky130_fd_sc_hd__nand2_2 _12631_ (.A(_03559_),
    .B(_03561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03562_));
 sky130_fd_sc_hd__o21ai_2 _12632_ (.A1(_03558_),
    .A2(_03560_),
    .B1(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03563_));
 sky130_fd_sc_hd__nor3_2 _12633_ (.A(_03535_),
    .B(_03558_),
    .C(_03560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03564_));
 sky130_fd_sc_hd__nand3b_2 _12634_ (.A_N(_03535_),
    .B(_03559_),
    .C(_03561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03565_));
 sky130_fd_sc_hd__nand2_2 _12635_ (.A(_03395_),
    .B(_03407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03566_));
 sky130_fd_sc_hd__a21oi_2 _12636_ (.A1(_03563_),
    .A2(_03565_),
    .B1(_03566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03567_));
 sky130_fd_sc_hd__a21o_2 _12637_ (.A1(_03563_),
    .A2(_03565_),
    .B1(_03566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03568_));
 sky130_fd_sc_hd__nand3_2 _12638_ (.A(_03563_),
    .B(_03565_),
    .C(_03566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03569_));
 sky130_fd_sc_hd__nand4_2 _12639_ (.A(_03532_),
    .B(_03533_),
    .C(_03568_),
    .D(_03569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03570_));
 sky130_fd_sc_hd__nand4_2 _12640_ (.A(_03395_),
    .B(_03407_),
    .C(_03563_),
    .D(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03571_));
 sky130_fd_sc_hd__a22o_2 _12641_ (.A1(_03395_),
    .A2(_03407_),
    .B1(_03563_),
    .B2(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03572_));
 sky130_fd_sc_hd__nand3_2 _12642_ (.A(_03534_),
    .B(_03571_),
    .C(_03572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03573_));
 sky130_fd_sc_hd__a21o_2 _12643_ (.A1(_03568_),
    .A2(_03569_),
    .B1(_03534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03574_));
 sky130_fd_sc_hd__nand3_2 _12644_ (.A(_03534_),
    .B(_03568_),
    .C(_03569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03575_));
 sky130_fd_sc_hd__nand3_2 _12645_ (.A(_03574_),
    .B(_03575_),
    .C(_03503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03576_));
 sky130_fd_sc_hd__and3_2 _12646_ (.A(_03504_),
    .B(_03570_),
    .C(_03573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03577_));
 sky130_fd_sc_hd__nand3_2 _12647_ (.A(_03504_),
    .B(_03570_),
    .C(_03573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_2 _12648_ (.A(_03576_),
    .B(_03578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03579_));
 sky130_fd_sc_hd__a41o_2 _12649_ (.A1(\a_h[6] ),
    .A2(\a_h[7] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_03402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03580_));
 sky130_fd_sc_hd__nand2_2 _12650_ (.A(_03412_),
    .B(_03413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03581_));
 sky130_fd_sc_hd__nand3_2 _12651_ (.A(_03411_),
    .B(_03580_),
    .C(_03581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03582_));
 sky130_fd_sc_hd__nand3b_2 _12652_ (.A_N(_03580_),
    .B(_03416_),
    .C(_03412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03583_));
 sky130_fd_sc_hd__nor2_2 _12653_ (.A(_09428_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03584_));
 sky130_fd_sc_hd__a21bo_2 _12654_ (.A1(_03582_),
    .A2(_03583_),
    .B1_N(_03584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03585_));
 sky130_fd_sc_hd__o211ai_2 _12655_ (.A1(_09428_),
    .A2(_09679_),
    .B1(_03582_),
    .C1(_03583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_2 _12656_ (.A(_03585_),
    .B(_03586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03587_));
 sky130_fd_sc_hd__a21oi_2 _12657_ (.A1(_03576_),
    .A2(_03578_),
    .B1(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03588_));
 sky130_fd_sc_hd__a21o_2 _12658_ (.A1(_03576_),
    .A2(_03578_),
    .B1(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03589_));
 sky130_fd_sc_hd__a32oi_2 _12659_ (.A1(_03574_),
    .A2(_03575_),
    .A3(_03503_),
    .B1(_03585_),
    .B2(_03586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03590_));
 sky130_fd_sc_hd__nand3_2 _12660_ (.A(_03576_),
    .B(_03578_),
    .C(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03591_));
 sky130_fd_sc_hd__nand4_2 _12661_ (.A(_03576_),
    .B(_03578_),
    .C(_03585_),
    .D(_03586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03592_));
 sky130_fd_sc_hd__nand2_2 _12662_ (.A(_03579_),
    .B(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03593_));
 sky130_fd_sc_hd__nand3_2 _12663_ (.A(_03593_),
    .B(_03501_),
    .C(_03592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03594_));
 sky130_fd_sc_hd__nand2_2 _12664_ (.A(_03502_),
    .B(_03591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03595_));
 sky130_fd_sc_hd__o21ai_2 _12665_ (.A1(_03588_),
    .A2(_03595_),
    .B1(_03594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_2 _12666_ (.A(_03596_),
    .B(_03500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03597_));
 sky130_fd_sc_hd__a31oi_2 _12667_ (.A1(_03593_),
    .A2(_03501_),
    .A3(_03592_),
    .B1(_03500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03598_));
 sky130_fd_sc_hd__o21ai_2 _12668_ (.A1(_03588_),
    .A2(_03595_),
    .B1(_03598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03599_));
 sky130_fd_sc_hd__a21o_2 _12669_ (.A1(_03597_),
    .A2(_03599_),
    .B1(_03499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03600_));
 sky130_fd_sc_hd__nand4b_2 _12670_ (.A_N(_03486_),
    .B(_03489_),
    .C(_03597_),
    .D(_03599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_2 _12671_ (.A(_03600_),
    .B(_03601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03602_));
 sky130_fd_sc_hd__nor2_2 _12672_ (.A(_03372_),
    .B(_03496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03603_));
 sky130_fd_sc_hd__o2111a_2 _12673_ (.A1(_03244_),
    .A2(_03248_),
    .B1(_03247_),
    .C1(_03114_),
    .D1(_03115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03604_));
 sky130_fd_sc_hd__nand4_2 _12674_ (.A(_03121_),
    .B(_03603_),
    .C(_03604_),
    .D(_03117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03605_));
 sky130_fd_sc_hd__o21ai_2 _12675_ (.A1(_03491_),
    .A2(_03370_),
    .B1(_03494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03606_));
 sky130_fd_sc_hd__a41oi_2 _12676_ (.A1(_03371_),
    .A2(_03373_),
    .A3(_03495_),
    .A4(_03247_),
    .B1(_03606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03607_));
 sky130_fd_sc_hd__nand3_2 _12677_ (.A(_03602_),
    .B(_03605_),
    .C(_03607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03608_));
 sky130_fd_sc_hd__a21o_2 _12678_ (.A1(_03605_),
    .A2(_03607_),
    .B1(_03602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03609_));
 sky130_fd_sc_hd__and3_2 _12679_ (.A(_09690_),
    .B(_03608_),
    .C(_03609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00294_));
 sky130_fd_sc_hd__a32oi_2 _12680_ (.A1(_03502_),
    .A2(_03589_),
    .A3(_03591_),
    .B1(_03594_),
    .B2(_03500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03610_));
 sky130_fd_sc_hd__a32o_2 _12681_ (.A1(_03502_),
    .A2(_03589_),
    .A3(_03591_),
    .B1(_03594_),
    .B2(_03500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03611_));
 sky130_fd_sc_hd__a21bo_2 _12682_ (.A1(_03583_),
    .A2(_03584_),
    .B1_N(_03582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03612_));
 sky130_fd_sc_hd__a32oi_2 _12683_ (.A1(_03504_),
    .A2(_03570_),
    .A3(_03573_),
    .B1(_03576_),
    .B2(_03587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03613_));
 sky130_fd_sc_hd__nor2_2 _12684_ (.A(_09439_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03614_));
 sky130_fd_sc_hd__o21ai_2 _12685_ (.A1(_03397_),
    .A2(_03550_),
    .B1(_03554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03615_));
 sky130_fd_sc_hd__a22oi_2 _12686_ (.A1(_03395_),
    .A2(_03407_),
    .B1(_03562_),
    .B2(_03535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_2 _12687_ (.A(_03563_),
    .B(_03566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03617_));
 sky130_fd_sc_hd__nand3b_2 _12688_ (.A_N(_03615_),
    .B(_03617_),
    .C(_03565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03618_));
 sky130_fd_sc_hd__o211ai_2 _12689_ (.A1(_03566_),
    .A2(_03564_),
    .B1(_03563_),
    .C1(_03615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03619_));
 sky130_fd_sc_hd__o311a_2 _12690_ (.A1(_03564_),
    .A2(_03615_),
    .A3(_03616_),
    .B1(_03614_),
    .C1(_03619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03620_));
 sky130_fd_sc_hd__nand4_2 _12691_ (.A(_03618_),
    .B(_03619_),
    .C(\a_h[6] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03621_));
 sky130_fd_sc_hd__a21oi_2 _12692_ (.A1(_03618_),
    .A2(_03619_),
    .B1(_03614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03622_));
 sky130_fd_sc_hd__a22o_2 _12693_ (.A1(\a_h[6] ),
    .A2(\b_h[15] ),
    .B1(_03618_),
    .B2(_03619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03623_));
 sky130_fd_sc_hd__nand2_2 _12694_ (.A(_03621_),
    .B(_03623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_2 _12695_ (.A(\a_h[8] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_2 _12696_ (.A(\a_h[9] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03626_));
 sky130_fd_sc_hd__and4_2 _12697_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03627_));
 sky130_fd_sc_hd__nand4_2 _12698_ (.A(\a_h[8] ),
    .B(\a_h[9] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03628_));
 sky130_fd_sc_hd__nand2_2 _12699_ (.A(_03625_),
    .B(_03626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03629_));
 sky130_fd_sc_hd__and4_2 _12700_ (.A(_03629_),
    .B(\b_h[14] ),
    .C(\a_h[7] ),
    .D(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03630_));
 sky130_fd_sc_hd__nand4_2 _12701_ (.A(_03629_),
    .B(\b_h[14] ),
    .C(\a_h[7] ),
    .D(_03628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03631_));
 sky130_fd_sc_hd__o2bb2a_2 _12702_ (.A1_N(_03628_),
    .A2_N(_03629_),
    .B1(_09449_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03632_));
 sky130_fd_sc_hd__a22o_2 _12703_ (.A1(\a_h[7] ),
    .A2(\b_h[14] ),
    .B1(_03628_),
    .B2(_03629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03633_));
 sky130_fd_sc_hd__nand2_2 _12704_ (.A(_03631_),
    .B(_03633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03634_));
 sky130_fd_sc_hd__and2_2 _12705_ (.A(\a_h[10] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03635_));
 sky130_fd_sc_hd__nand2_2 _12706_ (.A(\a_h[10] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2_2 _12707_ (.A(\a_h[11] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2_2 _12708_ (.A(\a_h[12] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03638_));
 sky130_fd_sc_hd__nand3_2 _12709_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03639_));
 sky130_fd_sc_hd__nand4_2 _12710_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03640_));
 sky130_fd_sc_hd__a22oi_2 _12711_ (.A1(\a_h[12] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_2 _12712_ (.A(_03637_),
    .B(_03638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03642_));
 sky130_fd_sc_hd__o21ai_2 _12713_ (.A1(_09635_),
    .A2(_03639_),
    .B1(_03642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03643_));
 sky130_fd_sc_hd__o2bb2ai_2 _12714_ (.A1_N(_03640_),
    .A2_N(_03642_),
    .B1(_09482_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03644_));
 sky130_fd_sc_hd__o211ai_2 _12715_ (.A1(_09635_),
    .A2(_03639_),
    .B1(_03635_),
    .C1(_03642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03645_));
 sky130_fd_sc_hd__nand2_2 _12716_ (.A(_03643_),
    .B(_03635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03646_));
 sky130_fd_sc_hd__o221ai_2 _12717_ (.A1(_09482_),
    .A2(_09646_),
    .B1(_03639_),
    .B2(_09635_),
    .C1(_03642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03647_));
 sky130_fd_sc_hd__nand2_2 _12718_ (.A(_03536_),
    .B(_03539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03648_));
 sky130_fd_sc_hd__o21ai_2 _12719_ (.A1(_03536_),
    .A2(_03540_),
    .B1(_03539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_2 _12720_ (.A(_03541_),
    .B(_03648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03650_));
 sky130_fd_sc_hd__and3_2 _12721_ (.A(_03646_),
    .B(_03647_),
    .C(_03650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03651_));
 sky130_fd_sc_hd__nand3_2 _12722_ (.A(_03646_),
    .B(_03647_),
    .C(_03650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03652_));
 sky130_fd_sc_hd__nand3_2 _12723_ (.A(_03644_),
    .B(_03649_),
    .C(_03645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03653_));
 sky130_fd_sc_hd__inv_2 _12724_ (.A(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03654_));
 sky130_fd_sc_hd__nand2_2 _12725_ (.A(_03652_),
    .B(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03655_));
 sky130_fd_sc_hd__o211ai_2 _12726_ (.A1(_03630_),
    .A2(_03632_),
    .B1(_03652_),
    .C1(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03656_));
 sky130_fd_sc_hd__a21o_2 _12727_ (.A1(_03652_),
    .A2(_03653_),
    .B1(_03634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03657_));
 sky130_fd_sc_hd__nand4_2 _12728_ (.A(_03631_),
    .B(_03633_),
    .C(_03652_),
    .D(_03653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03658_));
 sky130_fd_sc_hd__o21ai_2 _12729_ (.A1(_03630_),
    .A2(_03632_),
    .B1(_03655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03659_));
 sky130_fd_sc_hd__nand3_2 _12730_ (.A(_03524_),
    .B(_03656_),
    .C(_03657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03660_));
 sky130_fd_sc_hd__and3_2 _12731_ (.A(_03659_),
    .B(_03523_),
    .C(_03658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03661_));
 sky130_fd_sc_hd__nand3_2 _12732_ (.A(_03659_),
    .B(_03523_),
    .C(_03658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03662_));
 sky130_fd_sc_hd__a31oi_2 _12733_ (.A1(_03549_),
    .A2(_03555_),
    .A3(_03556_),
    .B1(_03547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03663_));
 sky130_fd_sc_hd__a31o_2 _12734_ (.A1(_03549_),
    .A2(_03555_),
    .A3(_03556_),
    .B1(_03547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03664_));
 sky130_fd_sc_hd__a21oi_2 _12735_ (.A1(_03660_),
    .A2(_03662_),
    .B1(_03663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03665_));
 sky130_fd_sc_hd__a21o_2 _12736_ (.A1(_03660_),
    .A2(_03662_),
    .B1(_03663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03666_));
 sky130_fd_sc_hd__a31oi_2 _12737_ (.A1(_03524_),
    .A2(_03656_),
    .A3(_03657_),
    .B1(_03664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03667_));
 sky130_fd_sc_hd__a31o_2 _12738_ (.A1(_03524_),
    .A2(_03656_),
    .A3(_03657_),
    .B1(_03664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03668_));
 sky130_fd_sc_hd__and3_2 _12739_ (.A(_03660_),
    .B(_03662_),
    .C(_03663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03669_));
 sky130_fd_sc_hd__nand3_2 _12740_ (.A(_03660_),
    .B(_03662_),
    .C(_03663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03670_));
 sky130_fd_sc_hd__o21ai_2 _12741_ (.A1(_03430_),
    .A2(_03507_),
    .B1(_03511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03671_));
 sky130_fd_sc_hd__a22o_2 _12742_ (.A1(\a_h[15] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03672_));
 sky130_fd_sc_hd__nand4_2 _12743_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03673_));
 sky130_fd_sc_hd__a22o_2 _12744_ (.A1(\a_h[13] ),
    .A2(\b_h[8] ),
    .B1(_03672_),
    .B2(_03673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03674_));
 sky130_fd_sc_hd__nand4_2 _12745_ (.A(_03672_),
    .B(_03673_),
    .C(\a_h[13] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03675_));
 sky130_fd_sc_hd__a21o_2 _12746_ (.A1(_03674_),
    .A2(_03675_),
    .B1(_03671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03676_));
 sky130_fd_sc_hd__and3_2 _12747_ (.A(_03671_),
    .B(_03674_),
    .C(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03677_));
 sky130_fd_sc_hd__nand3_2 _12748_ (.A(_03671_),
    .B(_03674_),
    .C(_03675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03678_));
 sky130_fd_sc_hd__nand2_2 _12749_ (.A(_03676_),
    .B(_03678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_2 _12750_ (.A(_03528_),
    .B(_03679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03680_));
 sky130_fd_sc_hd__inv_2 _12751_ (.A(_03680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03681_));
 sky130_fd_sc_hd__nand3b_2 _12752_ (.A_N(_03679_),
    .B(_03522_),
    .C(_03527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_2 _12753_ (.A(_03680_),
    .B(_03682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03683_));
 sky130_fd_sc_hd__o211ai_2 _12754_ (.A1(_03661_),
    .A2(_03668_),
    .B1(_03682_),
    .C1(_03666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03684_));
 sky130_fd_sc_hd__o21ai_2 _12755_ (.A1(_03665_),
    .A2(_03669_),
    .B1(_03683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03685_));
 sky130_fd_sc_hd__o21ai_2 _12756_ (.A1(_03681_),
    .A2(_03684_),
    .B1(_03685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03686_));
 sky130_fd_sc_hd__nand2_2 _12757_ (.A(_03532_),
    .B(_03569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03687_));
 sky130_fd_sc_hd__o22a_2 _12758_ (.A1(_03452_),
    .A2(_03531_),
    .B1(_03567_),
    .B2(_03687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03688_));
 sky130_fd_sc_hd__o22ai_2 _12759_ (.A1(_03452_),
    .A2(_03531_),
    .B1(_03567_),
    .B2(_03687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_2 _12760_ (.A(_03686_),
    .B(_03688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03690_));
 sky130_fd_sc_hd__o211ai_2 _12761_ (.A1(_03681_),
    .A2(_03684_),
    .B1(_03685_),
    .C1(_03689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03691_));
 sky130_fd_sc_hd__o211ai_2 _12762_ (.A1(_03620_),
    .A2(_03622_),
    .B1(_03690_),
    .C1(_03691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03692_));
 sky130_fd_sc_hd__a21o_2 _12763_ (.A1(_03690_),
    .A2(_03691_),
    .B1(_03624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03693_));
 sky130_fd_sc_hd__nand4_2 _12764_ (.A(_03621_),
    .B(_03623_),
    .C(_03690_),
    .D(_03691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03694_));
 sky130_fd_sc_hd__a22o_2 _12765_ (.A1(_03621_),
    .A2(_03623_),
    .B1(_03690_),
    .B2(_03691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03695_));
 sky130_fd_sc_hd__o211ai_2 _12766_ (.A1(_03577_),
    .A2(_03590_),
    .B1(_03694_),
    .C1(_03695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_2 _12767_ (.A(_03693_),
    .B(_03613_),
    .C(_03692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03697_));
 sky130_fd_sc_hd__a21o_2 _12768_ (.A1(_03696_),
    .A2(_03697_),
    .B1(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03698_));
 sky130_fd_sc_hd__nand3_2 _12769_ (.A(_03696_),
    .B(_03697_),
    .C(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03699_));
 sky130_fd_sc_hd__a21bo_2 _12770_ (.A1(_03696_),
    .A2(_03697_),
    .B1_N(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03700_));
 sky130_fd_sc_hd__nand3b_2 _12771_ (.A_N(_03612_),
    .B(_03696_),
    .C(_03697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03701_));
 sky130_fd_sc_hd__nand3_2 _12772_ (.A(_03611_),
    .B(_03698_),
    .C(_03699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03702_));
 sky130_fd_sc_hd__nand3_2 _12773_ (.A(_03700_),
    .B(_03701_),
    .C(_03610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03703_));
 sky130_fd_sc_hd__and2_2 _12774_ (.A(_03702_),
    .B(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_2 _12775_ (.A(_03702_),
    .B(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03705_));
 sky130_fd_sc_hd__nand2_2 _12776_ (.A(_03600_),
    .B(_03609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03706_));
 sky130_fd_sc_hd__a31o_2 _12777_ (.A1(_03600_),
    .A2(_03609_),
    .A3(_03705_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03707_));
 sky130_fd_sc_hd__a21oi_2 _12778_ (.A1(_03704_),
    .A2(_03706_),
    .B1(_03707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_2 _12779_ (.A(_03697_),
    .B(_03612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03708_));
 sky130_fd_sc_hd__nand2_2 _12780_ (.A(_03696_),
    .B(_03708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03709_));
 sky130_fd_sc_hd__a21boi_2 _12781_ (.A1(_03612_),
    .A2(_03697_),
    .B1_N(_03696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03710_));
 sky130_fd_sc_hd__a21bo_2 _12782_ (.A1(_03614_),
    .A2(_03618_),
    .B1_N(_03619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03711_));
 sky130_fd_sc_hd__inv_2 _12783_ (.A(_03711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03712_));
 sky130_fd_sc_hd__o21ai_2 _12784_ (.A1(_03620_),
    .A2(_03622_),
    .B1(_03691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_2 _12785_ (.A(_03690_),
    .B(_03713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03714_));
 sky130_fd_sc_hd__a21boi_2 _12786_ (.A1(_03624_),
    .A2(_03691_),
    .B1_N(_03690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03715_));
 sky130_fd_sc_hd__nor2_2 _12787_ (.A(_09449_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03716_));
 sky130_fd_sc_hd__a31o_2 _12788_ (.A1(\a_h[7] ),
    .A2(_03629_),
    .A3(\b_h[14] ),
    .B1(_03627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03717_));
 sky130_fd_sc_hd__o22a_2 _12789_ (.A1(_03627_),
    .A2(_03630_),
    .B1(_03661_),
    .B2(_03667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03718_));
 sky130_fd_sc_hd__o21ai_2 _12790_ (.A1(_03661_),
    .A2(_03667_),
    .B1(_03717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03719_));
 sky130_fd_sc_hd__nand3b_2 _12791_ (.A_N(_03717_),
    .B(_03668_),
    .C(_03662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03720_));
 sky130_fd_sc_hd__a21oi_2 _12792_ (.A1(_03719_),
    .A2(_03720_),
    .B1(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03721_));
 sky130_fd_sc_hd__a22o_2 _12793_ (.A1(\a_h[7] ),
    .A2(\b_h[15] ),
    .B1(_03719_),
    .B2(_03720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03722_));
 sky130_fd_sc_hd__nand2_2 _12794_ (.A(_03720_),
    .B(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03723_));
 sky130_fd_sc_hd__and3_2 _12795_ (.A(_03719_),
    .B(_03720_),
    .C(_03716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03724_));
 sky130_fd_sc_hd__o21ai_2 _12796_ (.A1(_03718_),
    .A2(_03723_),
    .B1(_03722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03725_));
 sky130_fd_sc_hd__nand2_2 _12797_ (.A(_03670_),
    .B(_03680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03726_));
 sky130_fd_sc_hd__o22ai_2 _12798_ (.A1(_03528_),
    .A2(_03679_),
    .B1(_03665_),
    .B2(_03726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03727_));
 sky130_fd_sc_hd__and4_2 _12799_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[7] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03728_));
 sky130_fd_sc_hd__a22oi_2 _12800_ (.A1(\a_h[15] ),
    .A2(\b_h[7] ),
    .B1(\b_h[8] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03729_));
 sky130_fd_sc_hd__nand3_2 _12801_ (.A(_03672_),
    .B(\b_h[8] ),
    .C(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03730_));
 sky130_fd_sc_hd__a211oi_2 _12802_ (.A1(_03673_),
    .A2(_03730_),
    .B1(_03729_),
    .C1(_03728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03731_));
 sky130_fd_sc_hd__a211o_2 _12803_ (.A1(_03673_),
    .A2(_03730_),
    .B1(_03729_),
    .C1(_03728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03732_));
 sky130_fd_sc_hd__o211a_2 _12804_ (.A1(_03728_),
    .A2(_03729_),
    .B1(_03730_),
    .C1(_03673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03733_));
 sky130_fd_sc_hd__or2_2 _12805_ (.A(_03731_),
    .B(_03733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03734_));
 sky130_fd_sc_hd__inv_2 _12806_ (.A(_03734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03735_));
 sky130_fd_sc_hd__and4_2 _12807_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03736_));
 sky130_fd_sc_hd__a22oi_2 _12808_ (.A1(\a_h[10] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03737_));
 sky130_fd_sc_hd__a22o_2 _12809_ (.A1(\a_h[10] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03738_));
 sky130_fd_sc_hd__o2111a_2 _12810_ (.A1(_02278_),
    .A2(_02589_),
    .B1(\a_h[8] ),
    .C1(\b_h[14] ),
    .D1(_03738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03739_));
 sky130_fd_sc_hd__o22a_2 _12811_ (.A1(_09460_),
    .A2(_09668_),
    .B1(_03736_),
    .B2(_03737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03740_));
 sky130_fd_sc_hd__nor2_2 _12812_ (.A(_03739_),
    .B(_03740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03741_));
 sky130_fd_sc_hd__o21ai_2 _12813_ (.A1(_03636_),
    .A2(_03641_),
    .B1(_03640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03742_));
 sky130_fd_sc_hd__o22a_2 _12814_ (.A1(_09635_),
    .A2(_03639_),
    .B1(_03636_),
    .B2(_03641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03743_));
 sky130_fd_sc_hd__nand2_2 _12815_ (.A(\a_h[11] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_2 _12816_ (.A(\a_h[12] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2_2 _12817_ (.A(\a_h[13] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03746_));
 sky130_fd_sc_hd__a22oi_2 _12818_ (.A1(\a_h[13] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_2 _12819_ (.A(_03745_),
    .B(_03746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03748_));
 sky130_fd_sc_hd__nand4_2 _12820_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03749_));
 sky130_fd_sc_hd__a21o_2 _12821_ (.A1(_03748_),
    .A2(_03749_),
    .B1(_03744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03750_));
 sky130_fd_sc_hd__o211ai_2 _12822_ (.A1(_09493_),
    .A2(_09646_),
    .B1(_03748_),
    .C1(_03749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03751_));
 sky130_fd_sc_hd__nand4_2 _12823_ (.A(_03748_),
    .B(_03749_),
    .C(\a_h[11] ),
    .D(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03752_));
 sky130_fd_sc_hd__a22o_2 _12824_ (.A1(\a_h[11] ),
    .A2(\b_h[11] ),
    .B1(_03748_),
    .B2(_03749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03753_));
 sky130_fd_sc_hd__nand3_2 _12825_ (.A(_03753_),
    .B(_03742_),
    .C(_03752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03754_));
 sky130_fd_sc_hd__inv_2 _12826_ (.A(_03754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03755_));
 sky130_fd_sc_hd__nand3_2 _12827_ (.A(_03743_),
    .B(_03750_),
    .C(_03751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_2 _12828_ (.A(_03754_),
    .B(_03756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03757_));
 sky130_fd_sc_hd__o21ai_2 _12829_ (.A1(_03739_),
    .A2(_03740_),
    .B1(_03756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_2 _12830_ (.A(_03757_),
    .B(_03741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03759_));
 sky130_fd_sc_hd__nand3_2 _12831_ (.A(_03741_),
    .B(_03754_),
    .C(_03756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03760_));
 sky130_fd_sc_hd__o21ai_2 _12832_ (.A1(_03739_),
    .A2(_03740_),
    .B1(_03757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03761_));
 sky130_fd_sc_hd__nand3_2 _12833_ (.A(_03761_),
    .B(_03677_),
    .C(_03760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03762_));
 sky130_fd_sc_hd__o211ai_2 _12834_ (.A1(_03758_),
    .A2(_03755_),
    .B1(_03678_),
    .C1(_03759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03763_));
 sky130_fd_sc_hd__and3_2 _12835_ (.A(_03631_),
    .B(_03633_),
    .C(_03652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03764_));
 sky130_fd_sc_hd__a31o_2 _12836_ (.A1(_03631_),
    .A2(_03633_),
    .A3(_03652_),
    .B1(_03654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03765_));
 sky130_fd_sc_hd__o2bb2ai_2 _12837_ (.A1_N(_03762_),
    .A2_N(_03763_),
    .B1(_03764_),
    .B2(_03654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03766_));
 sky130_fd_sc_hd__o2111ai_2 _12838_ (.A1(_03634_),
    .A2(_03651_),
    .B1(_03653_),
    .C1(_03762_),
    .D1(_03763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03767_));
 sky130_fd_sc_hd__o21ai_2 _12839_ (.A1(_03654_),
    .A2(_03764_),
    .B1(_03763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03768_));
 sky130_fd_sc_hd__o211ai_2 _12840_ (.A1(_03654_),
    .A2(_03764_),
    .B1(_03763_),
    .C1(_03762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03769_));
 sky130_fd_sc_hd__a21o_2 _12841_ (.A1(_03762_),
    .A2(_03763_),
    .B1(_03765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03770_));
 sky130_fd_sc_hd__nand2_2 _12842_ (.A(_03769_),
    .B(_03770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03771_));
 sky130_fd_sc_hd__nand3_2 _12843_ (.A(_03770_),
    .B(_03735_),
    .C(_03769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03772_));
 sky130_fd_sc_hd__nand3_2 _12844_ (.A(_03734_),
    .B(_03766_),
    .C(_03767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03773_));
 sky130_fd_sc_hd__nand3_2 _12845_ (.A(_03727_),
    .B(_03772_),
    .C(_03773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03774_));
 sky130_fd_sc_hd__a21oi_2 _12846_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03775_));
 sky130_fd_sc_hd__a21o_2 _12847_ (.A1(_03772_),
    .A2(_03773_),
    .B1(_03727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03776_));
 sky130_fd_sc_hd__a21o_2 _12848_ (.A1(_03774_),
    .A2(_03776_),
    .B1(_03725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03777_));
 sky130_fd_sc_hd__o211ai_2 _12849_ (.A1(_03721_),
    .A2(_03724_),
    .B1(_03774_),
    .C1(_03776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03778_));
 sky130_fd_sc_hd__nand3b_2 _12850_ (.A_N(_03725_),
    .B(_03774_),
    .C(_03776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03779_));
 sky130_fd_sc_hd__a2bb2o_2 _12851_ (.A1_N(_03721_),
    .A2_N(_03724_),
    .B1(_03774_),
    .B2(_03776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03780_));
 sky130_fd_sc_hd__and3_2 _12852_ (.A(_03715_),
    .B(_03779_),
    .C(_03780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03781_));
 sky130_fd_sc_hd__nand3_2 _12853_ (.A(_03715_),
    .B(_03779_),
    .C(_03780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03782_));
 sky130_fd_sc_hd__nand3_2 _12854_ (.A(_03714_),
    .B(_03777_),
    .C(_03778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03783_));
 sky130_fd_sc_hd__a31o_2 _12855_ (.A1(_03714_),
    .A2(_03777_),
    .A3(_03778_),
    .B1(_03712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03784_));
 sky130_fd_sc_hd__a21o_2 _12856_ (.A1(_03782_),
    .A2(_03783_),
    .B1(_03711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03785_));
 sky130_fd_sc_hd__o211ai_2 _12857_ (.A1(_03781_),
    .A2(_03784_),
    .B1(_03785_),
    .C1(_03709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03786_));
 sky130_fd_sc_hd__nand3_2 _12858_ (.A(_03712_),
    .B(_03782_),
    .C(_03783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03787_));
 sky130_fd_sc_hd__a21o_2 _12859_ (.A1(_03782_),
    .A2(_03783_),
    .B1(_03712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03788_));
 sky130_fd_sc_hd__nand3_2 _12860_ (.A(_03710_),
    .B(_03787_),
    .C(_03788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03789_));
 sky130_fd_sc_hd__and2_2 _12861_ (.A(_03786_),
    .B(_03789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03790_));
 sky130_fd_sc_hd__a21boi_2 _12862_ (.A1(_03600_),
    .A2(_03702_),
    .B1_N(_03703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03791_));
 sky130_fd_sc_hd__or2_2 _12863_ (.A(_03602_),
    .B(_03705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03792_));
 sky130_fd_sc_hd__a21oi_2 _12864_ (.A1(_03605_),
    .A2(_03607_),
    .B1(_03792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03793_));
 sky130_fd_sc_hd__o21ai_2 _12865_ (.A1(_03791_),
    .A2(_03793_),
    .B1(_03790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03794_));
 sky130_fd_sc_hd__o31a_2 _12866_ (.A1(_03790_),
    .A2(_03791_),
    .A3(_03793_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03795_));
 sky130_fd_sc_hd__and2_2 _12867_ (.A(_03795_),
    .B(_03794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00296_));
 sky130_fd_sc_hd__o21ai_2 _12868_ (.A1(_03775_),
    .A2(_03725_),
    .B1(_03774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03796_));
 sky130_fd_sc_hd__nor2_2 _12869_ (.A(_03736_),
    .B(_03739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03797_));
 sky130_fd_sc_hd__a31o_2 _12870_ (.A1(_03761_),
    .A2(_03677_),
    .A3(_03760_),
    .B1(_03765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03798_));
 sky130_fd_sc_hd__o211ai_2 _12871_ (.A1(_03736_),
    .A2(_03739_),
    .B1(_03763_),
    .C1(_03798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03799_));
 sky130_fd_sc_hd__nand3_2 _12872_ (.A(_03762_),
    .B(_03768_),
    .C(_03797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03800_));
 sky130_fd_sc_hd__nand2_2 _12873_ (.A(\a_h[8] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03801_));
 sky130_fd_sc_hd__o211ai_2 _12874_ (.A1(_09460_),
    .A2(_09679_),
    .B1(_03799_),
    .C1(_03800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03802_));
 sky130_fd_sc_hd__a21o_2 _12875_ (.A1(_03799_),
    .A2(_03800_),
    .B1(_03801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03803_));
 sky130_fd_sc_hd__a22o_2 _12876_ (.A1(\a_h[8] ),
    .A2(\b_h[15] ),
    .B1(_03799_),
    .B2(_03800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03804_));
 sky130_fd_sc_hd__nand4_2 _12877_ (.A(_03799_),
    .B(_03800_),
    .C(\a_h[8] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_2 _12878_ (.A(_03507_),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03806_));
 sky130_fd_sc_hd__and3_2 _12879_ (.A(_03507_),
    .B(\b_h[8] ),
    .C(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03807_));
 sky130_fd_sc_hd__a21o_2 _12880_ (.A1(_03741_),
    .A2(_03756_),
    .B1(_03755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03808_));
 sky130_fd_sc_hd__a21boi_2 _12881_ (.A1(_03741_),
    .A2(_03756_),
    .B1_N(_03754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2_2 _12882_ (.A(\a_h[10] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_2 _12883_ (.A(\a_h[11] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_2 _12884_ (.A(_03810_),
    .B(_03811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03812_));
 sky130_fd_sc_hd__nand4_2 _12885_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03813_));
 sky130_fd_sc_hd__and4_2 _12886_ (.A(_03812_),
    .B(_03813_),
    .C(\a_h[9] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03814_));
 sky130_fd_sc_hd__o2111ai_2 _12887_ (.A1(_02362_),
    .A2(_02589_),
    .B1(\a_h[9] ),
    .C1(\b_h[14] ),
    .D1(_03812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03815_));
 sky130_fd_sc_hd__o2bb2a_2 _12888_ (.A1_N(_03812_),
    .A2_N(_03813_),
    .B1(_09471_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03816_));
 sky130_fd_sc_hd__a22o_2 _12889_ (.A1(\a_h[9] ),
    .A2(\b_h[14] ),
    .B1(_03812_),
    .B2(_03813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03817_));
 sky130_fd_sc_hd__nor2_2 _12890_ (.A(_03814_),
    .B(_03816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03818_));
 sky130_fd_sc_hd__nand2_2 _12891_ (.A(_03815_),
    .B(_03817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03819_));
 sky130_fd_sc_hd__a21o_2 _12892_ (.A1(_03744_),
    .A2(_03749_),
    .B1(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03820_));
 sky130_fd_sc_hd__a21oi_2 _12893_ (.A1(_03744_),
    .A2(_03749_),
    .B1(_03747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03821_));
 sky130_fd_sc_hd__nor2_2 _12894_ (.A(_09504_),
    .B(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_2 _12895_ (.A(\a_h[12] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_2 _12896_ (.A(\a_h[13] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_2 _12897_ (.A(\a_h[14] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03825_));
 sky130_fd_sc_hd__nand3_2 _12898_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03826_));
 sky130_fd_sc_hd__and4_2 _12899_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03827_));
 sky130_fd_sc_hd__nand4_2 _12900_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_2 _12901_ (.A(_03824_),
    .B(_03825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03829_));
 sky130_fd_sc_hd__o21ai_2 _12902_ (.A1(_09635_),
    .A2(_03826_),
    .B1(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_2 _12903_ (.A(_03830_),
    .B(_03822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03831_));
 sky130_fd_sc_hd__o221ai_2 _12904_ (.A1(_09504_),
    .A2(_09646_),
    .B1(_03826_),
    .B2(_09635_),
    .C1(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03832_));
 sky130_fd_sc_hd__o2bb2ai_2 _12905_ (.A1_N(_03828_),
    .A2_N(_03829_),
    .B1(_09504_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03833_));
 sky130_fd_sc_hd__o2111ai_2 _12906_ (.A1(_09635_),
    .A2(_03826_),
    .B1(\b_h[11] ),
    .C1(\a_h[12] ),
    .D1(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03834_));
 sky130_fd_sc_hd__a21oi_2 _12907_ (.A1(_03833_),
    .A2(_03834_),
    .B1(_03821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03835_));
 sky130_fd_sc_hd__nand3_2 _12908_ (.A(_03831_),
    .B(_03832_),
    .C(_03820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03836_));
 sky130_fd_sc_hd__nand3_2 _12909_ (.A(_03821_),
    .B(_03833_),
    .C(_03834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_2 _12910_ (.A(_03836_),
    .B(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_2 _12911_ (.A(_03838_),
    .B(_03818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03839_));
 sky130_fd_sc_hd__o211ai_2 _12912_ (.A1(_03814_),
    .A2(_03816_),
    .B1(_03836_),
    .C1(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03840_));
 sky130_fd_sc_hd__nand4_2 _12913_ (.A(_03815_),
    .B(_03817_),
    .C(_03836_),
    .D(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03841_));
 sky130_fd_sc_hd__a22o_2 _12914_ (.A1(_03815_),
    .A2(_03817_),
    .B1(_03836_),
    .B2(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03842_));
 sky130_fd_sc_hd__a21oi_2 _12915_ (.A1(_03839_),
    .A2(_03840_),
    .B1(_03732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03843_));
 sky130_fd_sc_hd__nand3_2 _12916_ (.A(_03842_),
    .B(_03731_),
    .C(_03841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03844_));
 sky130_fd_sc_hd__nand3_2 _12917_ (.A(_03732_),
    .B(_03839_),
    .C(_03840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_2 _12918_ (.A(_03844_),
    .B(_03845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03846_));
 sky130_fd_sc_hd__a21oi_2 _12919_ (.A1(_03844_),
    .A2(_03845_),
    .B1(_03808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03847_));
 sky130_fd_sc_hd__a21o_2 _12920_ (.A1(_03844_),
    .A2(_03845_),
    .B1(_03808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03848_));
 sky130_fd_sc_hd__a31oi_2 _12921_ (.A1(_03732_),
    .A2(_03839_),
    .A3(_03840_),
    .B1(_03809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03849_));
 sky130_fd_sc_hd__a31o_2 _12922_ (.A1(_03732_),
    .A2(_03839_),
    .A3(_03840_),
    .B1(_03809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03850_));
 sky130_fd_sc_hd__nand2_2 _12923_ (.A(_03849_),
    .B(_03844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03851_));
 sky130_fd_sc_hd__a21oi_2 _12924_ (.A1(_03844_),
    .A2(_03849_),
    .B1(_03847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03852_));
 sky130_fd_sc_hd__nand3_2 _12925_ (.A(_03809_),
    .B(_03844_),
    .C(_03845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2_2 _12926_ (.A(_03846_),
    .B(_03808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03854_));
 sky130_fd_sc_hd__o211ai_2 _12927_ (.A1(_09613_),
    .A2(_03806_),
    .B1(_03853_),
    .C1(_03854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03855_));
 sky130_fd_sc_hd__nand3_2 _12928_ (.A(_03848_),
    .B(_03851_),
    .C(_03807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03856_));
 sky130_fd_sc_hd__nand3b_2 _12929_ (.A_N(_03772_),
    .B(_03855_),
    .C(_03856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03857_));
 sky130_fd_sc_hd__o2bb2ai_2 _12930_ (.A1_N(_03855_),
    .A2_N(_03856_),
    .B1(_03734_),
    .B2(_03771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03858_));
 sky130_fd_sc_hd__nand4_2 _12931_ (.A(_03802_),
    .B(_03803_),
    .C(_03857_),
    .D(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03859_));
 sky130_fd_sc_hd__a22o_2 _12932_ (.A1(_03802_),
    .A2(_03803_),
    .B1(_03857_),
    .B2(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03860_));
 sky130_fd_sc_hd__o2111a_2 _12933_ (.A1(_03775_),
    .A2(_03725_),
    .B1(_03774_),
    .C1(_03859_),
    .D1(_03860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03861_));
 sky130_fd_sc_hd__o2111ai_2 _12934_ (.A1(_03775_),
    .A2(_03725_),
    .B1(_03774_),
    .C1(_03859_),
    .D1(_03860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03862_));
 sky130_fd_sc_hd__nand3_2 _12935_ (.A(_03804_),
    .B(_03805_),
    .C(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03863_));
 sky130_fd_sc_hd__nand4_2 _12936_ (.A(_03804_),
    .B(_03805_),
    .C(_03857_),
    .D(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03864_));
 sky130_fd_sc_hd__a22o_2 _12937_ (.A1(_03804_),
    .A2(_03805_),
    .B1(_03857_),
    .B2(_03858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03865_));
 sky130_fd_sc_hd__nand3_2 _12938_ (.A(_03865_),
    .B(_03796_),
    .C(_03864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03866_));
 sky130_fd_sc_hd__and2_2 _12939_ (.A(_03862_),
    .B(_03866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03867_));
 sky130_fd_sc_hd__a31o_2 _12940_ (.A1(\a_h[7] ),
    .A2(_03720_),
    .A3(\b_h[15] ),
    .B1(_03718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03868_));
 sky130_fd_sc_hd__a21oi_2 _12941_ (.A1(_03862_),
    .A2(_03866_),
    .B1(_03868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03869_));
 sky130_fd_sc_hd__and3_2 _12942_ (.A(_03862_),
    .B(_03866_),
    .C(_03868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03870_));
 sky130_fd_sc_hd__a21boi_2 _12943_ (.A1(_03711_),
    .A2(_03783_),
    .B1_N(_03782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03871_));
 sky130_fd_sc_hd__o211a_2 _12944_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_03782_),
    .C1(_03784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03872_));
 sky130_fd_sc_hd__o21ai_2 _12945_ (.A1(_03869_),
    .A2(_03870_),
    .B1(_03871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03873_));
 sky130_fd_sc_hd__o2bb2ai_2 _12946_ (.A1_N(_03782_),
    .A2_N(_03784_),
    .B1(_03868_),
    .B2(_03867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03874_));
 sky130_fd_sc_hd__o21a_2 _12947_ (.A1(_03870_),
    .A2(_03874_),
    .B1(_03873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03875_));
 sky130_fd_sc_hd__nand2_2 _12948_ (.A(_03786_),
    .B(_03794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03876_));
 sky130_fd_sc_hd__o21ai_2 _12949_ (.A1(_03875_),
    .A2(_03876_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03877_));
 sky130_fd_sc_hd__a21oi_2 _12950_ (.A1(_03875_),
    .A2(_03876_),
    .B1(_03877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00297_));
 sky130_fd_sc_hd__a31o_2 _12951_ (.A1(_03719_),
    .A2(_03723_),
    .A3(_03866_),
    .B1(_03861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_2 _12952_ (.A(\a_h[9] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03879_));
 sky130_fd_sc_hd__a31o_2 _12953_ (.A1(\a_h[10] ),
    .A2(\a_h[11] ),
    .A3(_02588_),
    .B1(_03814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03880_));
 sky130_fd_sc_hd__o21ai_2 _12954_ (.A1(_03843_),
    .A2(_03849_),
    .B1(_03880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03881_));
 sky130_fd_sc_hd__nand3b_2 _12955_ (.A_N(_03880_),
    .B(_03850_),
    .C(_03844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_2 _12956_ (.A(_03881_),
    .B(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03883_));
 sky130_fd_sc_hd__nand4_2 _12957_ (.A(_03881_),
    .B(_03882_),
    .C(\a_h[9] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03884_));
 sky130_fd_sc_hd__a22o_2 _12958_ (.A1(\a_h[9] ),
    .A2(\b_h[15] ),
    .B1(_03881_),
    .B2(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03885_));
 sky130_fd_sc_hd__a21oi_2 _12959_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03886_));
 sky130_fd_sc_hd__a21o_2 _12960_ (.A1(_03881_),
    .A2(_03882_),
    .B1(_03879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03887_));
 sky130_fd_sc_hd__o211a_2 _12961_ (.A1(_09471_),
    .A2(_09679_),
    .B1(_03881_),
    .C1(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03888_));
 sky130_fd_sc_hd__o211ai_2 _12962_ (.A1(_09471_),
    .A2(_09679_),
    .B1(_03881_),
    .C1(_03882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03889_));
 sky130_fd_sc_hd__and2_2 _12963_ (.A(\a_h[10] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03890_));
 sky130_fd_sc_hd__nand2_2 _12964_ (.A(\a_h[12] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03891_));
 sky130_fd_sc_hd__nand4_2 _12965_ (.A(\a_h[11] ),
    .B(\a_h[12] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_2 _12966_ (.A(\a_h[11] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_2 _12967_ (.A(\a_h[12] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_2 _12968_ (.A(_03893_),
    .B(_03894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03895_));
 sky130_fd_sc_hd__and3_2 _12969_ (.A(_03895_),
    .B(_03890_),
    .C(_03892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03896_));
 sky130_fd_sc_hd__o2111ai_2 _12970_ (.A1(_02502_),
    .A2(_02589_),
    .B1(\a_h[10] ),
    .C1(\b_h[14] ),
    .D1(_03895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03897_));
 sky130_fd_sc_hd__a21oi_2 _12971_ (.A1(_03892_),
    .A2(_03895_),
    .B1(_03890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03898_));
 sky130_fd_sc_hd__a22o_2 _12972_ (.A1(\a_h[10] ),
    .A2(\b_h[14] ),
    .B1(_03892_),
    .B2(_03895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03899_));
 sky130_fd_sc_hd__nor2_2 _12973_ (.A(_03896_),
    .B(_03898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_2 _12974_ (.A(_03897_),
    .B(_03899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_2 _12975_ (.A(\a_h[13] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03902_));
 sky130_fd_sc_hd__and2_2 _12976_ (.A(\a_h[14] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03903_));
 sky130_fd_sc_hd__nand2_2 _12977_ (.A(\a_h[14] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03904_));
 sky130_fd_sc_hd__nand2_2 _12978_ (.A(\a_h[15] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03905_));
 sky130_fd_sc_hd__nand4_2 _12979_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03906_));
 sky130_fd_sc_hd__a22oi_2 _12980_ (.A1(\a_h[15] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03907_));
 sky130_fd_sc_hd__nand2_2 _12981_ (.A(_03904_),
    .B(_03905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03908_));
 sky130_fd_sc_hd__o2bb2ai_2 _12982_ (.A1_N(_03906_),
    .A2_N(_03908_),
    .B1(_09515_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03909_));
 sky130_fd_sc_hd__nand4_2 _12983_ (.A(_03908_),
    .B(\b_h[11] ),
    .C(\a_h[13] ),
    .D(_03906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03910_));
 sky130_fd_sc_hd__a21oi_2 _12984_ (.A1(_03824_),
    .A2(_03825_),
    .B1(_03823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03911_));
 sky130_fd_sc_hd__a21boi_2 _12985_ (.A1(_03823_),
    .A2(_03828_),
    .B1_N(_03829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03912_));
 sky130_fd_sc_hd__a21oi_2 _12986_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03913_));
 sky130_fd_sc_hd__a21o_2 _12987_ (.A1(_03909_),
    .A2(_03910_),
    .B1(_03912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03914_));
 sky130_fd_sc_hd__o211a_2 _12988_ (.A1(_03827_),
    .A2(_03911_),
    .B1(_03910_),
    .C1(_03909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03915_));
 sky130_fd_sc_hd__o2111ai_2 _12989_ (.A1(_03822_),
    .A2(_03827_),
    .B1(_03829_),
    .C1(_03909_),
    .D1(_03910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03916_));
 sky130_fd_sc_hd__nand3_2 _12990_ (.A(_03914_),
    .B(_03916_),
    .C(_03900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03917_));
 sky130_fd_sc_hd__o22ai_2 _12991_ (.A1(_03896_),
    .A2(_03898_),
    .B1(_03913_),
    .B2(_03915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03918_));
 sky130_fd_sc_hd__o21ai_2 _12992_ (.A1(_03913_),
    .A2(_03915_),
    .B1(_03900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03919_));
 sky130_fd_sc_hd__o211ai_2 _12993_ (.A1(_03896_),
    .A2(_03898_),
    .B1(_03914_),
    .C1(_03916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03920_));
 sky130_fd_sc_hd__nand3_2 _12994_ (.A(_03918_),
    .B(_03728_),
    .C(_03917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03921_));
 sky130_fd_sc_hd__a21oi_2 _12995_ (.A1(_03917_),
    .A2(_03918_),
    .B1(_03728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03922_));
 sky130_fd_sc_hd__nand3b_2 _12996_ (.A_N(_03728_),
    .B(_03919_),
    .C(_03920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03923_));
 sky130_fd_sc_hd__o21ai_2 _12997_ (.A1(_03819_),
    .A2(_03835_),
    .B1(_03837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03924_));
 sky130_fd_sc_hd__nand3_2 _12998_ (.A(_03921_),
    .B(_03923_),
    .C(_03924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03925_));
 sky130_fd_sc_hd__a21o_2 _12999_ (.A1(_03921_),
    .A2(_03923_),
    .B1(_03924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03926_));
 sky130_fd_sc_hd__nand2_2 _13000_ (.A(_03925_),
    .B(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03927_));
 sky130_fd_sc_hd__nor2_2 _13001_ (.A(_03856_),
    .B(_03927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03928_));
 sky130_fd_sc_hd__nand4_2 _13002_ (.A(_03807_),
    .B(_03852_),
    .C(_03925_),
    .D(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03929_));
 sky130_fd_sc_hd__a32oi_2 _13003_ (.A1(_03848_),
    .A2(_03851_),
    .A3(_03807_),
    .B1(_03925_),
    .B2(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03930_));
 sky130_fd_sc_hd__a32o_2 _13004_ (.A1(_03848_),
    .A2(_03851_),
    .A3(_03807_),
    .B1(_03925_),
    .B2(_03926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03931_));
 sky130_fd_sc_hd__o211ai_2 _13005_ (.A1(_03856_),
    .A2(_03927_),
    .B1(_03889_),
    .C1(_03887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03932_));
 sky130_fd_sc_hd__nand4_2 _13006_ (.A(_03887_),
    .B(_03889_),
    .C(_03929_),
    .D(_03931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03933_));
 sky130_fd_sc_hd__o22ai_2 _13007_ (.A1(_03886_),
    .A2(_03888_),
    .B1(_03928_),
    .B2(_03930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03934_));
 sky130_fd_sc_hd__nand4_2 _13008_ (.A(_03884_),
    .B(_03885_),
    .C(_03929_),
    .D(_03931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03935_));
 sky130_fd_sc_hd__o2bb2ai_2 _13009_ (.A1_N(_03884_),
    .A2_N(_03885_),
    .B1(_03928_),
    .B2(_03930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03936_));
 sky130_fd_sc_hd__nand3_2 _13010_ (.A(_03802_),
    .B(_03803_),
    .C(_03857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03937_));
 sky130_fd_sc_hd__nand4_2 _13011_ (.A(_03858_),
    .B(_03935_),
    .C(_03936_),
    .D(_03937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03938_));
 sky130_fd_sc_hd__nand4_2 _13012_ (.A(_03857_),
    .B(_03863_),
    .C(_03933_),
    .D(_03934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03939_));
 sky130_fd_sc_hd__nand2_2 _13013_ (.A(_03938_),
    .B(_03939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03940_));
 sky130_fd_sc_hd__a31o_2 _13014_ (.A1(_03762_),
    .A2(_03768_),
    .A3(_03797_),
    .B1(_03801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03941_));
 sky130_fd_sc_hd__nand2_2 _13015_ (.A(_03799_),
    .B(_03941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03942_));
 sky130_fd_sc_hd__inv_2 _13016_ (.A(_03942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03943_));
 sky130_fd_sc_hd__and3_2 _13017_ (.A(_03938_),
    .B(_03939_),
    .C(_03943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03944_));
 sky130_fd_sc_hd__or2_2 _13018_ (.A(_03942_),
    .B(_03940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03945_));
 sky130_fd_sc_hd__a22o_2 _13019_ (.A1(_03938_),
    .A2(_03939_),
    .B1(_03941_),
    .B2(_03799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03946_));
 sky130_fd_sc_hd__nand2_2 _13020_ (.A(_03878_),
    .B(_03946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03947_));
 sky130_fd_sc_hd__a21o_2 _13021_ (.A1(_03945_),
    .A2(_03946_),
    .B1(_03878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03948_));
 sky130_fd_sc_hd__o21a_2 _13022_ (.A1(_03944_),
    .A2(_03947_),
    .B1(_03948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03949_));
 sky130_fd_sc_hd__nand4_2 _13023_ (.A(_03791_),
    .B(_03875_),
    .C(_03786_),
    .D(_03789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03950_));
 sky130_fd_sc_hd__o32a_2 _13024_ (.A1(_03869_),
    .A2(_03870_),
    .A3(_03871_),
    .B1(_03786_),
    .B2(_03872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03951_));
 sky130_fd_sc_hd__nand4b_2 _13025_ (.A_N(_03602_),
    .B(_03704_),
    .C(_03790_),
    .D(_03875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03952_));
 sky130_fd_sc_hd__nand4_2 _13026_ (.A(_03605_),
    .B(_03607_),
    .C(_03950_),
    .D(_03951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03953_));
 sky130_fd_sc_hd__nand3_2 _13027_ (.A(_03950_),
    .B(_03952_),
    .C(_03951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03954_));
 sky130_fd_sc_hd__a21o_2 _13028_ (.A1(_03953_),
    .A2(_03954_),
    .B1(_03949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03955_));
 sky130_fd_sc_hd__o2111ai_2 _13029_ (.A1(_03944_),
    .A2(_03947_),
    .B1(_03948_),
    .C1(_03953_),
    .D1(_03954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03956_));
 sky130_fd_sc_hd__and3_2 _13030_ (.A(_09690_),
    .B(_03955_),
    .C(_03956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00298_));
 sky130_fd_sc_hd__o31a_2 _13031_ (.A1(_09471_),
    .A2(_09679_),
    .A3(_03883_),
    .B1(_03881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03957_));
 sky130_fd_sc_hd__o21ai_2 _13032_ (.A1(_03901_),
    .A2(_03913_),
    .B1(_03916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_2 _13033_ (.A(\a_h[13] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03959_));
 sky130_fd_sc_hd__nand4_2 _13034_ (.A(\a_h[12] ),
    .B(\a_h[13] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_2 _13035_ (.A(_03891_),
    .B(_03959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03961_));
 sky130_fd_sc_hd__o2bb2ai_2 _13036_ (.A1_N(_03960_),
    .A2_N(_03961_),
    .B1(_09493_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03962_));
 sky130_fd_sc_hd__nand4_2 _13037_ (.A(_03961_),
    .B(\b_h[14] ),
    .C(\a_h[11] ),
    .D(_03960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03963_));
 sky130_fd_sc_hd__and2_2 _13038_ (.A(\a_h[15] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03964_));
 sky130_fd_sc_hd__and4_2 _13039_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[10] ),
    .D(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03965_));
 sky130_fd_sc_hd__nand2_2 _13040_ (.A(_03903_),
    .B(_03964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03966_));
 sky130_fd_sc_hd__a22oi_2 _13041_ (.A1(\a_h[15] ),
    .A2(\b_h[10] ),
    .B1(\b_h[11] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03967_));
 sky130_fd_sc_hd__a21oi_2 _13042_ (.A1(_03903_),
    .A2(_03964_),
    .B1(_03967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03968_));
 sky130_fd_sc_hd__o21ai_2 _13043_ (.A1(_03902_),
    .A2(_03907_),
    .B1(_03906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03969_));
 sky130_fd_sc_hd__o221ai_2 _13044_ (.A1(_03904_),
    .A2(_03905_),
    .B1(_03965_),
    .B2(_03967_),
    .C1(_03910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_2 _13045_ (.A(_03969_),
    .B(_03968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03971_));
 sky130_fd_sc_hd__a22o_2 _13046_ (.A1(_03962_),
    .A2(_03963_),
    .B1(_03970_),
    .B2(_03971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03972_));
 sky130_fd_sc_hd__nand4_2 _13047_ (.A(_03962_),
    .B(_03963_),
    .C(_03970_),
    .D(_03971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_2 _13048_ (.A(_03972_),
    .B(_03973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03974_));
 sky130_fd_sc_hd__nand3_2 _13049_ (.A(_03958_),
    .B(_03972_),
    .C(_03973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03975_));
 sky130_fd_sc_hd__xnor2_2 _13050_ (.A(_03958_),
    .B(_03974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03976_));
 sky130_fd_sc_hd__nor2_2 _13051_ (.A(_09482_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03977_));
 sky130_fd_sc_hd__a31o_2 _13052_ (.A1(\a_h[11] ),
    .A2(\a_h[12] ),
    .A3(_02588_),
    .B1(_03896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03978_));
 sky130_fd_sc_hd__a31oi_2 _13053_ (.A1(_03918_),
    .A2(_03728_),
    .A3(_03917_),
    .B1(_03924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03979_));
 sky130_fd_sc_hd__a31o_2 _13054_ (.A1(_03918_),
    .A2(_03728_),
    .A3(_03917_),
    .B1(_03924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03980_));
 sky130_fd_sc_hd__o21bai_2 _13055_ (.A1(_03922_),
    .A2(_03979_),
    .B1_N(_03978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03981_));
 sky130_fd_sc_hd__nand3_2 _13056_ (.A(_03923_),
    .B(_03978_),
    .C(_03980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03982_));
 sky130_fd_sc_hd__nand4_2 _13057_ (.A(_03981_),
    .B(_03982_),
    .C(\a_h[10] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03983_));
 sky130_fd_sc_hd__a21o_2 _13058_ (.A1(_03981_),
    .A2(_03982_),
    .B1(_03977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03984_));
 sky130_fd_sc_hd__a31o_2 _13059_ (.A1(_03923_),
    .A2(_03978_),
    .A3(_03980_),
    .B1(_03977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03985_));
 sky130_fd_sc_hd__a21o_2 _13060_ (.A1(_03983_),
    .A2(_03984_),
    .B1(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03986_));
 sky130_fd_sc_hd__nand3_2 _13061_ (.A(_03984_),
    .B(_03976_),
    .C(_03983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03987_));
 sky130_fd_sc_hd__a22o_2 _13062_ (.A1(_03931_),
    .A2(_03932_),
    .B1(_03986_),
    .B2(_03987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03988_));
 sky130_fd_sc_hd__nand4_2 _13063_ (.A(_03931_),
    .B(_03932_),
    .C(_03986_),
    .D(_03987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03989_));
 sky130_fd_sc_hd__nand3b_2 _13064_ (.A_N(_03957_),
    .B(_03988_),
    .C(_03989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03990_));
 sky130_fd_sc_hd__a21bo_2 _13065_ (.A1(_03988_),
    .A2(_03989_),
    .B1_N(_03957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03991_));
 sky130_fd_sc_hd__o21ai_2 _13066_ (.A1(_03940_),
    .A2(_03943_),
    .B1(_03938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03992_));
 sky130_fd_sc_hd__a21oi_2 _13067_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03993_));
 sky130_fd_sc_hd__a21o_2 _13068_ (.A1(_03990_),
    .A2(_03991_),
    .B1(_03992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_03994_));
 sky130_fd_sc_hd__nand3_2 _13069_ (.A(_03990_),
    .B(_03991_),
    .C(_03992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_2 _13070_ (.A(_03994_),
    .B(_03995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03996_));
 sky130_fd_sc_hd__inv_2 _13071_ (.A(_03996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_2 _13072_ (.A(_03948_),
    .B(_03956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03998_));
 sky130_fd_sc_hd__a21oi_2 _13073_ (.A1(_03998_),
    .A2(_03997_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_03999_));
 sky130_fd_sc_hd__o21a_2 _13074_ (.A1(_03997_),
    .A2(_03998_),
    .B1(_03999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00299_));
 sky130_fd_sc_hd__and3_2 _13075_ (.A(_03904_),
    .B(\b_h[11] ),
    .C(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04000_));
 sky130_fd_sc_hd__nor2_2 _13076_ (.A(_09504_),
    .B(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_2 _13077_ (.A(\a_h[14] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04002_));
 sky130_fd_sc_hd__nand4_2 _13078_ (.A(\a_h[13] ),
    .B(\a_h[14] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04003_));
 sky130_fd_sc_hd__a22o_2 _13079_ (.A1(\a_h[14] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04004_));
 sky130_fd_sc_hd__o311a_2 _13080_ (.A1(_09515_),
    .A2(_09657_),
    .A3(_04002_),
    .B1(_04004_),
    .C1(_04001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04005_));
 sky130_fd_sc_hd__o2111ai_2 _13081_ (.A1(_03959_),
    .A2(_04002_),
    .B1(\a_h[12] ),
    .C1(\b_h[14] ),
    .D1(_04004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04006_));
 sky130_fd_sc_hd__a21oi_2 _13082_ (.A1(_04003_),
    .A2(_04004_),
    .B1(_04001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04007_));
 sky130_fd_sc_hd__o2bb2ai_2 _13083_ (.A1_N(_03964_),
    .A2_N(_03904_),
    .B1(_04007_),
    .B2(_04005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04008_));
 sky130_fd_sc_hd__nand3b_2 _13084_ (.A_N(_04007_),
    .B(_04000_),
    .C(_04006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04009_));
 sky130_fd_sc_hd__a22o_2 _13085_ (.A1(_03969_),
    .A2(_03968_),
    .B1(_03963_),
    .B2(_03962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04010_));
 sky130_fd_sc_hd__o21ai_2 _13086_ (.A1(_03968_),
    .A2(_03969_),
    .B1(_04010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04011_));
 sky130_fd_sc_hd__a22o_2 _13087_ (.A1(_04008_),
    .A2(_04009_),
    .B1(_04010_),
    .B2(_03970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04012_));
 sky130_fd_sc_hd__o2111ai_2 _13088_ (.A1(_03969_),
    .A2(_03968_),
    .B1(_04009_),
    .C1(_04008_),
    .D1(_04010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_2 _13089_ (.A(_04012_),
    .B(_04013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04014_));
 sky130_fd_sc_hd__o31a_2 _13090_ (.A1(_09515_),
    .A2(_09657_),
    .A3(_03891_),
    .B1(_03963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04015_));
 sky130_fd_sc_hd__o21ai_2 _13091_ (.A1(_03891_),
    .A2(_03959_),
    .B1(_03963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04016_));
 sky130_fd_sc_hd__nand4_2 _13092_ (.A(_03958_),
    .B(_03972_),
    .C(_03973_),
    .D(_04016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04017_));
 sky130_fd_sc_hd__nand2_2 _13093_ (.A(_03975_),
    .B(_04015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04018_));
 sky130_fd_sc_hd__o2bb2ai_2 _13094_ (.A1_N(_04017_),
    .A2_N(_04018_),
    .B1(_09493_),
    .B2(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04019_));
 sky130_fd_sc_hd__nand4_2 _13095_ (.A(_04018_),
    .B(\b_h[15] ),
    .C(\a_h[11] ),
    .D(_04017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04020_));
 sky130_fd_sc_hd__a22oi_2 _13096_ (.A1(_04012_),
    .A2(_04013_),
    .B1(_04019_),
    .B2(_04020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04021_));
 sky130_fd_sc_hd__a41oi_2 _13097_ (.A1(_04018_),
    .A2(\b_h[15] ),
    .A3(\a_h[11] ),
    .A4(_04017_),
    .B1(_04014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04022_));
 sky130_fd_sc_hd__a21oi_2 _13098_ (.A1(_04019_),
    .A2(_04022_),
    .B1(_04021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04023_));
 sky130_fd_sc_hd__nand4_2 _13099_ (.A(_03983_),
    .B(_04023_),
    .C(_03984_),
    .D(_03976_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04024_));
 sky130_fd_sc_hd__a31o_2 _13100_ (.A1(_03976_),
    .A2(_03983_),
    .A3(_03984_),
    .B1(_04023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04025_));
 sky130_fd_sc_hd__a22o_2 _13101_ (.A1(_03981_),
    .A2(_03985_),
    .B1(_04024_),
    .B2(_04025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04026_));
 sky130_fd_sc_hd__nand3_2 _13102_ (.A(_03981_),
    .B(_03985_),
    .C(_04025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04027_));
 sky130_fd_sc_hd__nand4_2 _13103_ (.A(_03981_),
    .B(_03985_),
    .C(_04024_),
    .D(_04025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2_2 _13104_ (.A(_03989_),
    .B(_03957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04029_));
 sky130_fd_sc_hd__a22o_2 _13105_ (.A1(_04026_),
    .A2(_04028_),
    .B1(_04029_),
    .B2(_03988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04030_));
 sky130_fd_sc_hd__and4_2 _13106_ (.A(_03988_),
    .B(_04026_),
    .C(_04028_),
    .D(_04029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04031_));
 sky130_fd_sc_hd__nand4_2 _13107_ (.A(_03988_),
    .B(_04026_),
    .C(_04028_),
    .D(_04029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04032_));
 sky130_fd_sc_hd__nand2_2 _13108_ (.A(_04030_),
    .B(_04032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04033_));
 sky130_fd_sc_hd__nand2_2 _13109_ (.A(_03949_),
    .B(_03997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04034_));
 sky130_fd_sc_hd__a31oi_2 _13110_ (.A1(_03950_),
    .A2(_03952_),
    .A3(_03951_),
    .B1(_04034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_2 _13111_ (.A(_03953_),
    .B(_04035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04036_));
 sky130_fd_sc_hd__o21a_2 _13112_ (.A1(_03993_),
    .A2(_03948_),
    .B1(_03995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04037_));
 sky130_fd_sc_hd__a21boi_2 _13113_ (.A1(_03953_),
    .A2(_04035_),
    .B1_N(_04037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04038_));
 sky130_fd_sc_hd__a21oi_2 _13114_ (.A1(_04036_),
    .A2(_04037_),
    .B1(_04033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04039_));
 sky130_fd_sc_hd__o21ai_2 _13115_ (.A1(_04033_),
    .A2(_04038_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04040_));
 sky130_fd_sc_hd__a21oi_2 _13116_ (.A1(_04033_),
    .A2(_04038_),
    .B1(_04040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00300_));
 sky130_fd_sc_hd__and4_2 _13117_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04041_));
 sky130_fd_sc_hd__nand4_2 _13118_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04042_));
 sky130_fd_sc_hd__a22o_2 _13119_ (.A1(\a_h[15] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04043_));
 sky130_fd_sc_hd__nand4_2 _13120_ (.A(_04043_),
    .B(\b_h[14] ),
    .C(\a_h[13] ),
    .D(_04042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04044_));
 sky130_fd_sc_hd__a22o_2 _13121_ (.A1(\a_h[13] ),
    .A2(\b_h[14] ),
    .B1(_04042_),
    .B2(_04043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04045_));
 sky130_fd_sc_hd__nand2_2 _13122_ (.A(_04044_),
    .B(_04045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04046_));
 sky130_fd_sc_hd__a21oi_2 _13123_ (.A1(_03966_),
    .A2(_04009_),
    .B1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04047_));
 sky130_fd_sc_hd__and3_2 _13124_ (.A(_03966_),
    .B(_04009_),
    .C(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04048_));
 sky130_fd_sc_hd__or2_2 _13125_ (.A(_04047_),
    .B(_04048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04049_));
 sky130_fd_sc_hd__o31a_2 _13126_ (.A1(_09515_),
    .A2(_09657_),
    .A3(_04002_),
    .B1(_04006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04050_));
 sky130_fd_sc_hd__a41o_2 _13127_ (.A1(\a_h[13] ),
    .A2(\a_h[14] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_04005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04051_));
 sky130_fd_sc_hd__and4b_2 _13128_ (.A_N(_04011_),
    .B(_04051_),
    .C(_04008_),
    .D(_04009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04052_));
 sky130_fd_sc_hd__nand4b_2 _13129_ (.A_N(_04011_),
    .B(_04051_),
    .C(_04008_),
    .D(_04009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_2 _13130_ (.A(_04013_),
    .B(_04050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04054_));
 sky130_fd_sc_hd__a211o_2 _13131_ (.A1(_04053_),
    .A2(_04054_),
    .B1(_09504_),
    .C1(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04055_));
 sky130_fd_sc_hd__o211ai_2 _13132_ (.A1(_09504_),
    .A2(_09679_),
    .B1(_04053_),
    .C1(_04054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04056_));
 sky130_fd_sc_hd__nand3_2 _13133_ (.A(_04049_),
    .B(_04055_),
    .C(_04056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04057_));
 sky130_fd_sc_hd__a21o_2 _13134_ (.A1(_04055_),
    .A2(_04056_),
    .B1(_04049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04058_));
 sky130_fd_sc_hd__nand4_2 _13135_ (.A(_04019_),
    .B(_04058_),
    .C(_04022_),
    .D(_04057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04059_));
 sky130_fd_sc_hd__a311o_2 _13136_ (.A1(_03960_),
    .A2(_03963_),
    .A3(_03975_),
    .B1(_09679_),
    .C1(_09493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04060_));
 sky130_fd_sc_hd__a22oi_2 _13137_ (.A1(_04022_),
    .A2(_04019_),
    .B1(_04058_),
    .B2(_04057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04061_));
 sky130_fd_sc_hd__a22o_2 _13138_ (.A1(_04022_),
    .A2(_04019_),
    .B1(_04058_),
    .B2(_04057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04062_));
 sky130_fd_sc_hd__a22o_2 _13139_ (.A1(_04017_),
    .A2(_04060_),
    .B1(_04062_),
    .B2(_04059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04063_));
 sky130_fd_sc_hd__nand4_2 _13140_ (.A(_04017_),
    .B(_04059_),
    .C(_04060_),
    .D(_04062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04064_));
 sky130_fd_sc_hd__a22oi_2 _13141_ (.A1(_04024_),
    .A2(_04027_),
    .B1(_04063_),
    .B2(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04065_));
 sky130_fd_sc_hd__nand4_2 _13142_ (.A(_04024_),
    .B(_04027_),
    .C(_04063_),
    .D(_04064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2b_2 _13143_ (.A_N(_04065_),
    .B(_04066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04067_));
 sky130_fd_sc_hd__o21ai_2 _13144_ (.A1(_04033_),
    .A2(_04038_),
    .B1(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04068_));
 sky130_fd_sc_hd__o21bai_2 _13145_ (.A1(_04031_),
    .A2(_04039_),
    .B1_N(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04069_));
 sky130_fd_sc_hd__o211a_2 _13146_ (.A1(_04068_),
    .A2(_04031_),
    .B1(_09690_),
    .C1(_04069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00301_));
 sky130_fd_sc_hd__a31o_2 _13147_ (.A1(_04017_),
    .A2(_04059_),
    .A3(_04060_),
    .B1(_04061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04070_));
 sky130_fd_sc_hd__a31o_2 _13148_ (.A1(_04054_),
    .A2(\b_h[15] ),
    .A3(\a_h[12] ),
    .B1(_04052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04071_));
 sky130_fd_sc_hd__a311oi_2 _13149_ (.A1(\a_h[13] ),
    .A2(_04043_),
    .A3(\b_h[14] ),
    .B1(_04041_),
    .C1(_04047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04072_));
 sky130_fd_sc_hd__a221oi_2 _13150_ (.A1(_03966_),
    .A2(_04009_),
    .B1(_04042_),
    .B2(_04044_),
    .C1(_04046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04073_));
 sky130_fd_sc_hd__nor4_2 _13151_ (.A(_09515_),
    .B(_04073_),
    .C(_09679_),
    .D(_04072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04074_));
 sky130_fd_sc_hd__o22a_2 _13152_ (.A1(_09515_),
    .A2(_09679_),
    .B1(_04072_),
    .B2(_04073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04075_));
 sky130_fd_sc_hd__a22o_2 _13153_ (.A1(\a_h[15] ),
    .A2(\b_h[13] ),
    .B1(\b_h[14] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04076_));
 sky130_fd_sc_hd__nand4_2 _13154_ (.A(\a_h[14] ),
    .B(\a_h[15] ),
    .C(\b_h[13] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04077_));
 sky130_fd_sc_hd__and4bb_2 _13155_ (.A_N(_04074_),
    .B_N(_04075_),
    .C(_04076_),
    .D(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04078_));
 sky130_fd_sc_hd__a2bb2oi_2 _13156_ (.A1_N(_04074_),
    .A2_N(_04075_),
    .B1(_04076_),
    .B2(_04077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04079_));
 sky130_fd_sc_hd__o21ai_2 _13157_ (.A1(_04078_),
    .A2(_04079_),
    .B1(_04058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04080_));
 sky130_fd_sc_hd__nor3_2 _13158_ (.A(_04079_),
    .B(_04058_),
    .C(_04078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04081_));
 sky130_fd_sc_hd__inv_2 _13159_ (.A(_04081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04082_));
 sky130_fd_sc_hd__a21o_2 _13160_ (.A1(_04080_),
    .A2(_04082_),
    .B1(_04071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04083_));
 sky130_fd_sc_hd__nand2_2 _13161_ (.A(_04080_),
    .B(_04071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04084_));
 sky130_fd_sc_hd__o21ai_2 _13162_ (.A1(_04081_),
    .A2(_04084_),
    .B1(_04083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04085_));
 sky130_fd_sc_hd__or2_2 _13163_ (.A(_04070_),
    .B(_04085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04086_));
 sky130_fd_sc_hd__xnor2_2 _13164_ (.A(_04070_),
    .B(_04085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04087_));
 sky130_fd_sc_hd__o21ai_2 _13165_ (.A1(_04031_),
    .A2(_04065_),
    .B1(_04066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04088_));
 sky130_fd_sc_hd__nor2_2 _13166_ (.A(_04033_),
    .B(_04067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04089_));
 sky130_fd_sc_hd__o31ai_2 _13167_ (.A1(_04033_),
    .A2(_04037_),
    .A3(_04067_),
    .B1(_04088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04090_));
 sky130_fd_sc_hd__o2111ai_2 _13168_ (.A1(_03944_),
    .A2(_03947_),
    .B1(_04089_),
    .C1(_03948_),
    .D1(_03997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04091_));
 sky130_fd_sc_hd__a31oi_2 _13169_ (.A1(_03950_),
    .A2(_03952_),
    .A3(_03951_),
    .B1(_04091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04092_));
 sky130_fd_sc_hd__a21o_2 _13170_ (.A1(_03953_),
    .A2(_04092_),
    .B1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04093_));
 sky130_fd_sc_hd__a21oi_2 _13171_ (.A1(_03953_),
    .A2(_04092_),
    .B1(_04090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04094_));
 sky130_fd_sc_hd__o21ai_2 _13172_ (.A1(_04087_),
    .A2(_04094_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_2 _13173_ (.A1(_04087_),
    .A2(_04094_),
    .B1(_04095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00302_));
 sky130_fd_sc_hd__or2_2 _13174_ (.A(_04073_),
    .B(_04074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_2 _13175_ (.A(\a_h[15] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_2 _13176_ (.A(\a_h[14] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04098_));
 sky130_fd_sc_hd__o22a_2 _13177_ (.A1(\b_h[15] ),
    .A2(_04002_),
    .B1(_04098_),
    .B2(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04099_));
 sky130_fd_sc_hd__or3b_2 _13178_ (.A(_04099_),
    .B(_09668_),
    .C_N(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04100_));
 sky130_fd_sc_hd__a22o_2 _13179_ (.A1(\a_h[15] ),
    .A2(\b_h[14] ),
    .B1(\b_h[15] ),
    .B2(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04101_));
 sky130_fd_sc_hd__a21o_2 _13180_ (.A1(_04100_),
    .A2(_04101_),
    .B1(_04078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04102_));
 sky130_fd_sc_hd__inv_2 _13181_ (.A(_04102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04103_));
 sky130_fd_sc_hd__and3_2 _13182_ (.A(_04078_),
    .B(_04100_),
    .C(_04101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04104_));
 sky130_fd_sc_hd__o21ai_2 _13183_ (.A1(_04103_),
    .A2(_04104_),
    .B1(_04096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04105_));
 sky130_fd_sc_hd__or3_2 _13184_ (.A(_04104_),
    .B(_04096_),
    .C(_04103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04106_));
 sky130_fd_sc_hd__nand2_2 _13185_ (.A(_04105_),
    .B(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04107_));
 sky130_fd_sc_hd__o21a_2 _13186_ (.A1(_04071_),
    .A2(_04081_),
    .B1(_04080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04108_));
 sky130_fd_sc_hd__a22o_2 _13187_ (.A1(_04082_),
    .A2(_04084_),
    .B1(_04105_),
    .B2(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04109_));
 sky130_fd_sc_hd__o311a_2 _13188_ (.A1(_04104_),
    .A2(_04096_),
    .A3(_04103_),
    .B1(_04084_),
    .C1(_04082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04110_));
 sky130_fd_sc_hd__and4_2 _13189_ (.A(_04082_),
    .B(_04084_),
    .C(_04105_),
    .D(_04106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04111_));
 sky130_fd_sc_hd__a21bo_2 _13190_ (.A1(_04105_),
    .A2(_04110_),
    .B1_N(_04109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04112_));
 sky130_fd_sc_hd__inv_2 _13191_ (.A(_04112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04113_));
 sky130_fd_sc_hd__o21ai_2 _13192_ (.A1(_04087_),
    .A2(_04094_),
    .B1(_04086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04114_));
 sky130_fd_sc_hd__o211ai_2 _13193_ (.A1(_04087_),
    .A2(_04094_),
    .B1(_04112_),
    .C1(_04086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04115_));
 sky130_fd_sc_hd__nand2_2 _13194_ (.A(_09690_),
    .B(_04115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04116_));
 sky130_fd_sc_hd__a21oi_2 _13195_ (.A1(_04113_),
    .A2(_04114_),
    .B1(_04116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00303_));
 sky130_fd_sc_hd__o2bb2a_2 _13196_ (.A1_N(\a_h[15] ),
    .A2_N(\b_h[15] ),
    .B1(_04097_),
    .B2(_04099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04117_));
 sky130_fd_sc_hd__a41o_2 _13197_ (.A1(\a_h[14] ),
    .A2(\a_h[15] ),
    .A3(\b_h[14] ),
    .A4(\b_h[15] ),
    .B1(_04117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04118_));
 sky130_fd_sc_hd__a21oi_2 _13198_ (.A1(_04096_),
    .A2(_04102_),
    .B1(_04104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04119_));
 sky130_fd_sc_hd__xnor2_2 _13199_ (.A(_04118_),
    .B(_04119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04120_));
 sky130_fd_sc_hd__inv_2 _13200_ (.A(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04121_));
 sky130_fd_sc_hd__o2bb2a_2 _13201_ (.A1_N(_04107_),
    .A2_N(_04108_),
    .B1(_04070_),
    .B2(_04085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04122_));
 sky130_fd_sc_hd__o31a_2 _13202_ (.A1(_04070_),
    .A2(_04085_),
    .A3(_04111_),
    .B1(_04109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04123_));
 sky130_fd_sc_hd__nor2_2 _13203_ (.A(_04087_),
    .B(_04112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04124_));
 sky130_fd_sc_hd__or3b_2 _13204_ (.A(_04111_),
    .B(_04087_),
    .C_N(_04109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04125_));
 sky130_fd_sc_hd__nand2_2 _13205_ (.A(_04093_),
    .B(_04124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04126_));
 sky130_fd_sc_hd__o21ai_2 _13206_ (.A1(_04094_),
    .A2(_04125_),
    .B1(_04123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04127_));
 sky130_fd_sc_hd__o221ai_2 _13207_ (.A1(_04111_),
    .A2(_04122_),
    .B1(_04125_),
    .B2(_04094_),
    .C1(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04128_));
 sky130_fd_sc_hd__a21oi_2 _13208_ (.A1(_04126_),
    .A2(_04123_),
    .B1(_04120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_2 _13209_ (.A(_04127_),
    .B(_04121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_2 _13210_ (.A(_09690_),
    .B(_04128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04131_));
 sky130_fd_sc_hd__nor2_2 _13211_ (.A(_04129_),
    .B(_04131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00304_));
 sky130_fd_sc_hd__o22a_2 _13212_ (.A1(_04097_),
    .A2(_04098_),
    .B1(_04117_),
    .B2(_04119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04132_));
 sky130_fd_sc_hd__a21oi_2 _13213_ (.A1(_04130_),
    .A2(_04132_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00305_));
 sky130_fd_sc_hd__and3_2 _13214_ (.A(_09690_),
    .B(\a_h[0] ),
    .C(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00306_));
 sky130_fd_sc_hd__and2_2 _13215_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04133_));
 sky130_fd_sc_hd__nand2_2 _13216_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04134_));
 sky130_fd_sc_hd__a22o_2 _13217_ (.A1(\b_l[1] ),
    .A2(\a_h[0] ),
    .B1(\a_h[1] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04135_));
 sky130_fd_sc_hd__o211a_2 _13218_ (.A1(_01855_),
    .A2(_04134_),
    .B1(_04135_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00307_));
 sky130_fd_sc_hd__and4_2 _13219_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04136_));
 sky130_fd_sc_hd__or2_2 _13220_ (.A(_01860_),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04137_));
 sky130_fd_sc_hd__a22o_2 _13221_ (.A1(\b_l[1] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04138_));
 sky130_fd_sc_hd__o2bb2a_2 _13222_ (.A1_N(_04137_),
    .A2_N(_04138_),
    .B1(_09155_),
    .B2(_09177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04139_));
 sky130_fd_sc_hd__and4_2 _13223_ (.A(_04138_),
    .B(\a_h[0] ),
    .C(\b_l[2] ),
    .D(_04137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_2 _13224_ (.A(_04139_),
    .B(_04140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04141_));
 sky130_fd_sc_hd__a31oi_2 _13225_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04133_),
    .B1(_04141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04142_));
 sky130_fd_sc_hd__and4_2 _13226_ (.A(_04141_),
    .B(_04133_),
    .C(\a_h[1] ),
    .D(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04143_));
 sky130_fd_sc_hd__nor3_2 _13227_ (.A(rst),
    .B(_04142_),
    .C(_04143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_2 _13228_ (.A(\a_h[0] ),
    .B(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04144_));
 sky130_fd_sc_hd__a31o_2 _13229_ (.A1(_04138_),
    .A2(\a_h[0] ),
    .A3(\b_l[2] ),
    .B1(_04136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04145_));
 sky130_fd_sc_hd__and4_2 _13230_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04146_));
 sky130_fd_sc_hd__nand4_2 _13231_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04147_));
 sky130_fd_sc_hd__a22o_2 _13232_ (.A1(\b_l[1] ),
    .A2(\a_h[2] ),
    .B1(\a_h[3] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04148_));
 sky130_fd_sc_hd__a22o_2 _13233_ (.A1(\b_l[2] ),
    .A2(\a_h[1] ),
    .B1(_04147_),
    .B2(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04149_));
 sky130_fd_sc_hd__o2111ai_2 _13234_ (.A1(_01871_),
    .A2(_04134_),
    .B1(\b_l[2] ),
    .C1(\a_h[1] ),
    .D1(_04148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04150_));
 sky130_fd_sc_hd__a21oi_2 _13235_ (.A1(_04149_),
    .A2(_04150_),
    .B1(_04145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04151_));
 sky130_fd_sc_hd__nand3_2 _13236_ (.A(_04145_),
    .B(_04149_),
    .C(_04150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2b_2 _13237_ (.A_N(_04151_),
    .B(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04153_));
 sky130_fd_sc_hd__xor2_2 _13238_ (.A(_04144_),
    .B(_04153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04154_));
 sky130_fd_sc_hd__a41o_2 _13239_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04133_),
    .A4(_04141_),
    .B1(_04154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04155_));
 sky130_fd_sc_hd__nand2_2 _13240_ (.A(_04143_),
    .B(_04154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04156_));
 sky130_fd_sc_hd__and3_2 _13241_ (.A(_09690_),
    .B(_04155_),
    .C(_04156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00309_));
 sky130_fd_sc_hd__and4_2 _13242_ (.A(\a_h[0] ),
    .B(\b_l[3] ),
    .C(\b_l[4] ),
    .D(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04157_));
 sky130_fd_sc_hd__a22oi_2 _13243_ (.A1(\a_h[0] ),
    .A2(\b_l[4] ),
    .B1(\a_h[1] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04158_));
 sky130_fd_sc_hd__or2_2 _13244_ (.A(_04157_),
    .B(_04158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04159_));
 sky130_fd_sc_hd__a31o_2 _13245_ (.A1(_04148_),
    .A2(\a_h[1] ),
    .A3(\b_l[2] ),
    .B1(_04146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04160_));
 sky130_fd_sc_hd__nand2_2 _13246_ (.A(\b_l[2] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_2 _13247_ (.A(\b_l[0] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04162_));
 sky130_fd_sc_hd__and4_2 _13248_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[3] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04163_));
 sky130_fd_sc_hd__nand4_2 _13249_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[3] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04164_));
 sky130_fd_sc_hd__a22oi_2 _13250_ (.A1(\b_l[1] ),
    .A2(\a_h[3] ),
    .B1(\a_h[4] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04165_));
 sky130_fd_sc_hd__o21ai_2 _13251_ (.A1(_04163_),
    .A2(_04165_),
    .B1(_04161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04166_));
 sky130_fd_sc_hd__nand4b_2 _13252_ (.A_N(_04165_),
    .B(\a_h[2] ),
    .C(\b_l[2] ),
    .D(_04164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04167_));
 sky130_fd_sc_hd__nand3_2 _13253_ (.A(_04160_),
    .B(_04166_),
    .C(_04167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04168_));
 sky130_fd_sc_hd__a21oi_2 _13254_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04169_));
 sky130_fd_sc_hd__a21o_2 _13255_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_04160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04170_));
 sky130_fd_sc_hd__a2bb2o_2 _13256_ (.A1_N(_04157_),
    .A2_N(_04158_),
    .B1(_04168_),
    .B2(_04170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04171_));
 sky130_fd_sc_hd__or4bb_2 _13257_ (.A(_04157_),
    .B(_04158_),
    .C_N(_04168_),
    .D_N(_04170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04172_));
 sky130_fd_sc_hd__o21ai_2 _13258_ (.A1(_04144_),
    .A2(_04151_),
    .B1(_04152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04173_));
 sky130_fd_sc_hd__nand3_2 _13259_ (.A(_04171_),
    .B(_04172_),
    .C(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04174_));
 sky130_fd_sc_hd__a21o_2 _13260_ (.A1(_04171_),
    .A2(_04172_),
    .B1(_04173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04175_));
 sky130_fd_sc_hd__nand2_2 _13261_ (.A(_04174_),
    .B(_04175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04176_));
 sky130_fd_sc_hd__a22o_2 _13262_ (.A1(_04143_),
    .A2(_04154_),
    .B1(_04174_),
    .B2(_04175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04177_));
 sky130_fd_sc_hd__or2_2 _13263_ (.A(_04156_),
    .B(_04176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04178_));
 sky130_fd_sc_hd__and3_2 _13264_ (.A(_09690_),
    .B(_04177_),
    .C(_04178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00310_));
 sky130_fd_sc_hd__o21ai_2 _13265_ (.A1(_04159_),
    .A2(_04169_),
    .B1(_04168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04179_));
 sky130_fd_sc_hd__o21a_2 _13266_ (.A1(_04159_),
    .A2(_04169_),
    .B1(_04168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04180_));
 sky130_fd_sc_hd__a22o_2 _13267_ (.A1(\b_l[4] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04181_));
 sky130_fd_sc_hd__nand2_2 _13268_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_2 _13269_ (.A(\b_l[4] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04183_));
 sky130_fd_sc_hd__and4_2 _13270_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04184_));
 sky130_fd_sc_hd__nand4_2 _13271_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04185_));
 sky130_fd_sc_hd__a22o_2 _13272_ (.A1(\a_h[0] ),
    .A2(\b_l[5] ),
    .B1(_04181_),
    .B2(_04185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04186_));
 sky130_fd_sc_hd__o211ai_2 _13273_ (.A1(_01860_),
    .A2(_04182_),
    .B1(\b_l[5] ),
    .C1(_04181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04187_));
 sky130_fd_sc_hd__and4_2 _13274_ (.A(_04181_),
    .B(_04185_),
    .C(\a_h[0] ),
    .D(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04188_));
 sky130_fd_sc_hd__o21ai_2 _13275_ (.A1(_09177_),
    .A2(_04187_),
    .B1(_04186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04189_));
 sky130_fd_sc_hd__nor2_2 _13276_ (.A(_04161_),
    .B(_04165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04190_));
 sky130_fd_sc_hd__o21ai_2 _13277_ (.A1(_04161_),
    .A2(_04165_),
    .B1(_04164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_2 _13278_ (.A(\b_l[2] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04192_));
 sky130_fd_sc_hd__a22oi_2 _13279_ (.A1(\b_l[1] ),
    .A2(\a_h[4] ),
    .B1(\a_h[5] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04193_));
 sky130_fd_sc_hd__a22o_2 _13280_ (.A1(\b_l[1] ),
    .A2(\a_h[4] ),
    .B1(\a_h[5] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04194_));
 sky130_fd_sc_hd__nand2_2 _13281_ (.A(\b_l[1] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04195_));
 sky130_fd_sc_hd__nor2_2 _13282_ (.A(_04162_),
    .B(_04195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04196_));
 sky130_fd_sc_hd__nand4_2 _13283_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04197_));
 sky130_fd_sc_hd__o21ai_2 _13284_ (.A1(_04193_),
    .A2(_04196_),
    .B1(_04192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04198_));
 sky130_fd_sc_hd__o2111ai_2 _13285_ (.A1(_04162_),
    .A2(_04195_),
    .B1(\b_l[2] ),
    .C1(\a_h[3] ),
    .D1(_04194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04199_));
 sky130_fd_sc_hd__a21o_2 _13286_ (.A1(_04198_),
    .A2(_04199_),
    .B1(_04191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04200_));
 sky130_fd_sc_hd__o211ai_2 _13287_ (.A1(_04163_),
    .A2(_04190_),
    .B1(_04198_),
    .C1(_04199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04201_));
 sky130_fd_sc_hd__a21o_2 _13288_ (.A1(_04200_),
    .A2(_04201_),
    .B1(_04189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04202_));
 sky130_fd_sc_hd__nand3_2 _13289_ (.A(_04189_),
    .B(_04200_),
    .C(_04201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04203_));
 sky130_fd_sc_hd__a21o_2 _13290_ (.A1(_04202_),
    .A2(_04203_),
    .B1(_04180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04204_));
 sky130_fd_sc_hd__nand3b_2 _13291_ (.A_N(_04179_),
    .B(_04202_),
    .C(_04203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04205_));
 sky130_fd_sc_hd__a21oi_2 _13292_ (.A1(_04204_),
    .A2(_04205_),
    .B1(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04206_));
 sky130_fd_sc_hd__and2_2 _13293_ (.A(_04205_),
    .B(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04207_));
 sky130_fd_sc_hd__nand2_2 _13294_ (.A(_04205_),
    .B(_04157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04208_));
 sky130_fd_sc_hd__a21o_2 _13295_ (.A1(_04207_),
    .A2(_04204_),
    .B1(_04206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04209_));
 sky130_fd_sc_hd__o21a_2 _13296_ (.A1(_04156_),
    .A2(_04176_),
    .B1(_04174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04210_));
 sky130_fd_sc_hd__a21o_2 _13297_ (.A1(_04174_),
    .A2(_04178_),
    .B1(_04209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_2 _13298_ (.A(_04210_),
    .B(_04209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04212_));
 sky130_fd_sc_hd__and3_2 _13299_ (.A(_04211_),
    .B(_04212_),
    .C(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00311_));
 sky130_fd_sc_hd__a211o_2 _13300_ (.A1(\a_h[0] ),
    .A2(\b_l[6] ),
    .B1(_04184_),
    .C1(_04188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04213_));
 sky130_fd_sc_hd__o211ai_2 _13301_ (.A1(_04184_),
    .A2(_04188_),
    .B1(\a_h[0] ),
    .C1(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04214_));
 sky130_fd_sc_hd__nand2_2 _13302_ (.A(_04213_),
    .B(_04214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_2 _13303_ (.A(_04189_),
    .B(_04201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04216_));
 sky130_fd_sc_hd__nand2_2 _13304_ (.A(_04200_),
    .B(_04216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04217_));
 sky130_fd_sc_hd__a21o_2 _13305_ (.A1(_04192_),
    .A2(_04197_),
    .B1(_04193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04218_));
 sky130_fd_sc_hd__a21oi_2 _13306_ (.A1(_04192_),
    .A2(_04197_),
    .B1(_04193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_2 _13307_ (.A(\b_l[2] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04220_));
 sky130_fd_sc_hd__nand2_2 _13308_ (.A(\b_l[1] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_2 _13309_ (.A(\b_l[0] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04222_));
 sky130_fd_sc_hd__nand4_2 _13310_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04223_));
 sky130_fd_sc_hd__a22oi_2 _13311_ (.A1(\b_l[1] ),
    .A2(\a_h[5] ),
    .B1(\a_h[6] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04224_));
 sky130_fd_sc_hd__nand2_2 _13312_ (.A(_04195_),
    .B(_04222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04225_));
 sky130_fd_sc_hd__o2bb2ai_2 _13313_ (.A1_N(_04223_),
    .A2_N(_04225_),
    .B1(_09155_),
    .B2(_09417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04226_));
 sky130_fd_sc_hd__nand4_2 _13314_ (.A(_04225_),
    .B(\a_h[4] ),
    .C(\b_l[2] ),
    .D(_04223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04227_));
 sky130_fd_sc_hd__o211ai_2 _13315_ (.A1(_09155_),
    .A2(_09417_),
    .B1(_04223_),
    .C1(_04225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04228_));
 sky130_fd_sc_hd__a21o_2 _13316_ (.A1(_04223_),
    .A2(_04225_),
    .B1(_04220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04229_));
 sky130_fd_sc_hd__a21oi_2 _13317_ (.A1(_04226_),
    .A2(_04227_),
    .B1(_04219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04230_));
 sky130_fd_sc_hd__nand3_2 _13318_ (.A(_04229_),
    .B(_04218_),
    .C(_04228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04231_));
 sky130_fd_sc_hd__nand3_2 _13319_ (.A(_04219_),
    .B(_04226_),
    .C(_04227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_2 _13320_ (.A(_04231_),
    .B(_04232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_2 _13321_ (.A(\b_l[5] ),
    .B(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_2 _13322_ (.A(\b_l[3] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04235_));
 sky130_fd_sc_hd__nand4_2 _13323_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04236_));
 sky130_fd_sc_hd__a22oi_2 _13324_ (.A1(\b_l[4] ),
    .A2(\a_h[2] ),
    .B1(\a_h[3] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_2 _13325_ (.A(_04183_),
    .B(_04235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04238_));
 sky130_fd_sc_hd__a22o_2 _13326_ (.A1(\b_l[5] ),
    .A2(\a_h[1] ),
    .B1(_04236_),
    .B2(_04238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04239_));
 sky130_fd_sc_hd__nand4_2 _13327_ (.A(_04238_),
    .B(\a_h[1] ),
    .C(\b_l[5] ),
    .D(_04236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_2 _13328_ (.A(_04239_),
    .B(_04240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_2 _13329_ (.A(_04233_),
    .B(_04241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04242_));
 sky130_fd_sc_hd__nand4_2 _13330_ (.A(_04231_),
    .B(_04232_),
    .C(_04239_),
    .D(_04240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_2 _13331_ (.A(_04242_),
    .B(_04243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04244_));
 sky130_fd_sc_hd__a22oi_2 _13332_ (.A1(_04200_),
    .A2(_04216_),
    .B1(_04242_),
    .B2(_04243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_2 _13333_ (.A(_04217_),
    .B(_04244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04246_));
 sky130_fd_sc_hd__nand4_2 _13334_ (.A(_04200_),
    .B(_04216_),
    .C(_04242_),
    .D(_04243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04247_));
 sky130_fd_sc_hd__a22o_2 _13335_ (.A1(_04213_),
    .A2(_04214_),
    .B1(_04246_),
    .B2(_04247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04248_));
 sky130_fd_sc_hd__nand4_2 _13336_ (.A(_04213_),
    .B(_04214_),
    .C(_04246_),
    .D(_04247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_2 _13337_ (.A(_04248_),
    .B(_04249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04250_));
 sky130_fd_sc_hd__inv_2 _13338_ (.A(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_2 _13339_ (.A(_04204_),
    .B(_04208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04252_));
 sky130_fd_sc_hd__a21o_2 _13340_ (.A1(_04248_),
    .A2(_04249_),
    .B1(_04252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04253_));
 sky130_fd_sc_hd__a21o_2 _13341_ (.A1(_04204_),
    .A2(_04208_),
    .B1(_04250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04254_));
 sky130_fd_sc_hd__nand2_2 _13342_ (.A(_04253_),
    .B(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04255_));
 sky130_fd_sc_hd__a21oi_2 _13343_ (.A1(_04211_),
    .A2(_04255_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04256_));
 sky130_fd_sc_hd__o31a_2 _13344_ (.A1(_04209_),
    .A2(_04210_),
    .A3(_04255_),
    .B1(_04256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00312_));
 sky130_fd_sc_hd__o21ai_2 _13345_ (.A1(_04215_),
    .A2(_04245_),
    .B1(_04247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04257_));
 sky130_fd_sc_hd__o21a_2 _13346_ (.A1(_04215_),
    .A2(_04245_),
    .B1(_04247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04258_));
 sky130_fd_sc_hd__and2_2 _13347_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04259_));
 sky130_fd_sc_hd__nand2_2 _13348_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04260_));
 sky130_fd_sc_hd__and3_2 _13349_ (.A(\a_h[0] ),
    .B(\a_h[1] ),
    .C(_04259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04261_));
 sky130_fd_sc_hd__a22oi_2 _13350_ (.A1(\a_h[0] ),
    .A2(\b_l[7] ),
    .B1(\a_h[1] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04262_));
 sky130_fd_sc_hd__a31o_2 _13351_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04259_),
    .B1(_04262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04263_));
 sky130_fd_sc_hd__a21o_2 _13352_ (.A1(_04234_),
    .A2(_04236_),
    .B1(_04237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04264_));
 sky130_fd_sc_hd__nor2_2 _13353_ (.A(_04264_),
    .B(_04263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04265_));
 sky130_fd_sc_hd__a311o_2 _13354_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04259_),
    .B1(_04262_),
    .C1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04266_));
 sky130_fd_sc_hd__o21ai_2 _13355_ (.A1(_04261_),
    .A2(_04262_),
    .B1(_04264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04267_));
 sky130_fd_sc_hd__and2_2 _13356_ (.A(_04266_),
    .B(_04267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04268_));
 sky130_fd_sc_hd__a21o_2 _13357_ (.A1(_04241_),
    .A2(_04232_),
    .B1(_04230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04269_));
 sky130_fd_sc_hd__a21oi_2 _13358_ (.A1(_04241_),
    .A2(_04232_),
    .B1(_04230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04270_));
 sky130_fd_sc_hd__nand2_2 _13359_ (.A(\b_l[5] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04271_));
 sky130_fd_sc_hd__nand4_2 _13360_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[3] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04272_));
 sky130_fd_sc_hd__a22oi_2 _13361_ (.A1(\b_l[4] ),
    .A2(\a_h[3] ),
    .B1(\a_h[4] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04273_));
 sky130_fd_sc_hd__a22o_2 _13362_ (.A1(\b_l[4] ),
    .A2(\a_h[3] ),
    .B1(\a_h[4] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04274_));
 sky130_fd_sc_hd__a22oi_2 _13363_ (.A1(\b_l[5] ),
    .A2(\a_h[2] ),
    .B1(_04272_),
    .B2(_04274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04275_));
 sky130_fd_sc_hd__and3_2 _13364_ (.A(_04272_),
    .B(\a_h[2] ),
    .C(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04276_));
 sky130_fd_sc_hd__and4_2 _13365_ (.A(_04274_),
    .B(\a_h[2] ),
    .C(\b_l[5] ),
    .D(_04272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04277_));
 sky130_fd_sc_hd__o221a_2 _13366_ (.A1(_09220_),
    .A2(_09395_),
    .B1(_01888_),
    .B2(_04182_),
    .C1(_04274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04278_));
 sky130_fd_sc_hd__a21oi_2 _13367_ (.A1(_04272_),
    .A2(_04274_),
    .B1(_04271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04279_));
 sky130_fd_sc_hd__a21oi_2 _13368_ (.A1(_04274_),
    .A2(_04276_),
    .B1(_04275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04280_));
 sky130_fd_sc_hd__a21o_2 _13369_ (.A1(_04220_),
    .A2(_04223_),
    .B1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04281_));
 sky130_fd_sc_hd__a21oi_2 _13370_ (.A1(_04220_),
    .A2(_04223_),
    .B1(_04224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04282_));
 sky130_fd_sc_hd__nand2_2 _13371_ (.A(\b_l[2] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_2 _13372_ (.A(\b_l[0] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04284_));
 sky130_fd_sc_hd__a22oi_2 _13373_ (.A1(\b_l[1] ),
    .A2(\a_h[6] ),
    .B1(\a_h[7] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_2 _13374_ (.A(_04221_),
    .B(_04284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04286_));
 sky130_fd_sc_hd__nand2_2 _13375_ (.A(\b_l[1] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04287_));
 sky130_fd_sc_hd__nand4_2 _13376_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[6] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04288_));
 sky130_fd_sc_hd__nand3_2 _13377_ (.A(_04288_),
    .B(\a_h[5] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04289_));
 sky130_fd_sc_hd__o2bb2ai_2 _13378_ (.A1_N(_04286_),
    .A2_N(_04288_),
    .B1(_09155_),
    .B2(_09428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04290_));
 sky130_fd_sc_hd__o221ai_2 _13379_ (.A1(_09155_),
    .A2(_09428_),
    .B1(_04222_),
    .B2(_04287_),
    .C1(_04286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04291_));
 sky130_fd_sc_hd__a21o_2 _13380_ (.A1(_04286_),
    .A2(_04288_),
    .B1(_04283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04292_));
 sky130_fd_sc_hd__o211a_2 _13381_ (.A1(_04289_),
    .A2(_04285_),
    .B1(_04282_),
    .C1(_04290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04293_));
 sky130_fd_sc_hd__o211ai_2 _13382_ (.A1(_04289_),
    .A2(_04285_),
    .B1(_04282_),
    .C1(_04290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04294_));
 sky130_fd_sc_hd__nand3_2 _13383_ (.A(_04292_),
    .B(_04281_),
    .C(_04291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_2 _13384_ (.A(_04294_),
    .B(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_2 _13385_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04297_));
 sky130_fd_sc_hd__o211ai_2 _13386_ (.A1(_04275_),
    .A2(_04277_),
    .B1(_04294_),
    .C1(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04298_));
 sky130_fd_sc_hd__o21ai_2 _13387_ (.A1(_04278_),
    .A2(_04279_),
    .B1(_04295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04299_));
 sky130_fd_sc_hd__a21o_2 _13388_ (.A1(_04294_),
    .A2(_04295_),
    .B1(_04280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04300_));
 sky130_fd_sc_hd__a21oi_2 _13389_ (.A1(_04297_),
    .A2(_04298_),
    .B1(_04269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04301_));
 sky130_fd_sc_hd__o211ai_2 _13390_ (.A1(_04299_),
    .A2(_04293_),
    .B1(_04270_),
    .C1(_04300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04302_));
 sky130_fd_sc_hd__nand3_2 _13391_ (.A(_04269_),
    .B(_04297_),
    .C(_04298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04303_));
 sky130_fd_sc_hd__nand3b_2 _13392_ (.A_N(_04268_),
    .B(_04302_),
    .C(_04303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04304_));
 sky130_fd_sc_hd__a21bo_2 _13393_ (.A1(_04302_),
    .A2(_04303_),
    .B1_N(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04305_));
 sky130_fd_sc_hd__a21o_2 _13394_ (.A1(_04302_),
    .A2(_04303_),
    .B1(_04268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04306_));
 sky130_fd_sc_hd__nand4_2 _13395_ (.A(_04266_),
    .B(_04267_),
    .C(_04302_),
    .D(_04303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04307_));
 sky130_fd_sc_hd__nand3_2 _13396_ (.A(_04258_),
    .B(_04304_),
    .C(_04305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04308_));
 sky130_fd_sc_hd__nand3_2 _13397_ (.A(_04306_),
    .B(_04307_),
    .C(_04257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04309_));
 sky130_fd_sc_hd__nand3_2 _13398_ (.A(_04214_),
    .B(_04308_),
    .C(_04309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04310_));
 sky130_fd_sc_hd__a21o_2 _13399_ (.A1(_04308_),
    .A2(_04309_),
    .B1(_04214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04311_));
 sky130_fd_sc_hd__nand2_2 _13400_ (.A(_04310_),
    .B(_04311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04312_));
 sky130_fd_sc_hd__nand3_2 _13401_ (.A(_04254_),
    .B(_04310_),
    .C(_04311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04313_));
 sky130_fd_sc_hd__a21o_2 _13402_ (.A1(_04310_),
    .A2(_04311_),
    .B1(_04254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04314_));
 sky130_fd_sc_hd__o2bb2a_2 _13403_ (.A1_N(_04313_),
    .A2_N(_04314_),
    .B1(_04255_),
    .B2(_04211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04315_));
 sky130_fd_sc_hd__nor3b_2 _13404_ (.A(_04174_),
    .B(_04209_),
    .C_N(_04253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_2 _13405_ (.A(_04316_),
    .B(_04313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04317_));
 sky130_fd_sc_hd__nor4b_2 _13406_ (.A(_04178_),
    .B(_04209_),
    .C(_04255_),
    .D_N(_04312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04318_));
 sky130_fd_sc_hd__a2111oi_2 _13407_ (.A1(_04313_),
    .A2(_04316_),
    .B1(_04318_),
    .C1(_04315_),
    .D1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00313_));
 sky130_fd_sc_hd__a21o_2 _13408_ (.A1(_04268_),
    .A2(_04303_),
    .B1(_04301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04319_));
 sky130_fd_sc_hd__a21oi_2 _13409_ (.A1(_04303_),
    .A2(_04268_),
    .B1(_04301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04320_));
 sky130_fd_sc_hd__nand4_2 _13410_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04321_));
 sky130_fd_sc_hd__a22o_2 _13411_ (.A1(\b_l[7] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04322_));
 sky130_fd_sc_hd__o2bb2ai_2 _13412_ (.A1_N(_04321_),
    .A2_N(_04322_),
    .B1(_09177_),
    .B2(_09264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04323_));
 sky130_fd_sc_hd__o2111ai_2 _13413_ (.A1(_01860_),
    .A2(_04260_),
    .B1(\a_h[0] ),
    .C1(\b_l[8] ),
    .D1(_04322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04324_));
 sky130_fd_sc_hd__a21oi_2 _13414_ (.A1(_04271_),
    .A2(_04272_),
    .B1(_04273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04325_));
 sky130_fd_sc_hd__a21oi_2 _13415_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04326_));
 sky130_fd_sc_hd__a21o_2 _13416_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04327_));
 sky130_fd_sc_hd__and3_2 _13417_ (.A(_04323_),
    .B(_04324_),
    .C(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04328_));
 sky130_fd_sc_hd__nand3_2 _13418_ (.A(_04323_),
    .B(_04324_),
    .C(_04325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04329_));
 sky130_fd_sc_hd__nand2_2 _13419_ (.A(_04327_),
    .B(_04261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04330_));
 sky130_fd_sc_hd__o211ai_2 _13420_ (.A1(_01855_),
    .A2(_04260_),
    .B1(_04327_),
    .C1(_04329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04331_));
 sky130_fd_sc_hd__o21ai_2 _13421_ (.A1(_04326_),
    .A2(_04328_),
    .B1(_04261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_2 _13422_ (.A(_04331_),
    .B(_04332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04333_));
 sky130_fd_sc_hd__nand2_2 _13423_ (.A(_04294_),
    .B(_04299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04334_));
 sky130_fd_sc_hd__a21oi_2 _13424_ (.A1(_04280_),
    .A2(_04295_),
    .B1(_04293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04335_));
 sky130_fd_sc_hd__nand2_2 _13425_ (.A(\b_l[5] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_2 _13426_ (.A(\b_l[4] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04337_));
 sky130_fd_sc_hd__nand4_2 _13427_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04338_));
 sky130_fd_sc_hd__nand2_2 _13428_ (.A(\b_l[4] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_2 _13429_ (.A(\b_l[3] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04340_));
 sky130_fd_sc_hd__a22oi_2 _13430_ (.A1(\b_l[4] ),
    .A2(\a_h[4] ),
    .B1(\a_h[5] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04341_));
 sky130_fd_sc_hd__nand2_2 _13431_ (.A(_04339_),
    .B(_04340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04342_));
 sky130_fd_sc_hd__o211ai_2 _13432_ (.A1(_09220_),
    .A2(_09406_),
    .B1(_04338_),
    .C1(_04342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04343_));
 sky130_fd_sc_hd__a21o_2 _13433_ (.A1(_04338_),
    .A2(_04342_),
    .B1(_04336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04344_));
 sky130_fd_sc_hd__nand2_2 _13434_ (.A(_04343_),
    .B(_04344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04345_));
 sky130_fd_sc_hd__a21o_2 _13435_ (.A1(_04283_),
    .A2(_04288_),
    .B1(_04285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04346_));
 sky130_fd_sc_hd__a21oi_2 _13436_ (.A1(_04283_),
    .A2(_04288_),
    .B1(_04285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2_2 _13437_ (.A(\b_l[2] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04348_));
 sky130_fd_sc_hd__nand2_2 _13438_ (.A(\b_l[0] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04349_));
 sky130_fd_sc_hd__a22oi_2 _13439_ (.A1(\b_l[1] ),
    .A2(\a_h[7] ),
    .B1(\a_h[8] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04350_));
 sky130_fd_sc_hd__nand2_2 _13440_ (.A(_04287_),
    .B(_04349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04351_));
 sky130_fd_sc_hd__nand4_2 _13441_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04352_));
 sky130_fd_sc_hd__a22oi_2 _13442_ (.A1(\b_l[2] ),
    .A2(\a_h[6] ),
    .B1(_04351_),
    .B2(_04352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04353_));
 sky130_fd_sc_hd__a41o_2 _13443_ (.A1(\b_l[0] ),
    .A2(\b_l[1] ),
    .A3(\a_h[7] ),
    .A4(\a_h[8] ),
    .B1(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04354_));
 sky130_fd_sc_hd__a21o_2 _13444_ (.A1(_04351_),
    .A2(_04352_),
    .B1(_04348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04355_));
 sky130_fd_sc_hd__o221ai_2 _13445_ (.A1(_09155_),
    .A2(_09439_),
    .B1(_02082_),
    .B2(_04134_),
    .C1(_04351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04356_));
 sky130_fd_sc_hd__o21ai_2 _13446_ (.A1(_04350_),
    .A2(_04354_),
    .B1(_04347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04357_));
 sky130_fd_sc_hd__nand3_2 _13447_ (.A(_04355_),
    .B(_04356_),
    .C(_04346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04358_));
 sky130_fd_sc_hd__o21ai_2 _13448_ (.A1(_04353_),
    .A2(_04357_),
    .B1(_04358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04359_));
 sky130_fd_sc_hd__o211ai_2 _13449_ (.A1(_04353_),
    .A2(_04357_),
    .B1(_04358_),
    .C1(_04345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04360_));
 sky130_fd_sc_hd__nand3_2 _13450_ (.A(_04343_),
    .B(_04344_),
    .C(_04359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04361_));
 sky130_fd_sc_hd__o2111ai_2 _13451_ (.A1(_04353_),
    .A2(_04357_),
    .B1(_04358_),
    .C1(_04344_),
    .D1(_04343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04362_));
 sky130_fd_sc_hd__nand2_2 _13452_ (.A(_04359_),
    .B(_04345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04363_));
 sky130_fd_sc_hd__a21oi_2 _13453_ (.A1(_04362_),
    .A2(_04363_),
    .B1(_04335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04364_));
 sky130_fd_sc_hd__nand3_2 _13454_ (.A(_04361_),
    .B(_04334_),
    .C(_04360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04365_));
 sky130_fd_sc_hd__nand3_2 _13455_ (.A(_04335_),
    .B(_04362_),
    .C(_04363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_2 _13456_ (.A(_04365_),
    .B(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04367_));
 sky130_fd_sc_hd__nand4_2 _13457_ (.A(_04331_),
    .B(_04332_),
    .C(_04365_),
    .D(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_2 _13458_ (.A(_04367_),
    .B(_04333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04369_));
 sky130_fd_sc_hd__nand3_2 _13459_ (.A(_04333_),
    .B(_04365_),
    .C(_04366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04370_));
 sky130_fd_sc_hd__a21o_2 _13460_ (.A1(_04365_),
    .A2(_04366_),
    .B1(_04333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04371_));
 sky130_fd_sc_hd__nand3_2 _13461_ (.A(_04371_),
    .B(_04319_),
    .C(_04370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04372_));
 sky130_fd_sc_hd__and3_2 _13462_ (.A(_04320_),
    .B(_04368_),
    .C(_04369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04373_));
 sky130_fd_sc_hd__nand3_2 _13463_ (.A(_04320_),
    .B(_04368_),
    .C(_04369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04374_));
 sky130_fd_sc_hd__a21o_2 _13464_ (.A1(_04372_),
    .A2(_04374_),
    .B1(_04265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04375_));
 sky130_fd_sc_hd__nand3_2 _13465_ (.A(_04372_),
    .B(_04374_),
    .C(_04265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04376_));
 sky130_fd_sc_hd__o211ai_2 _13466_ (.A1(_04264_),
    .A2(_04263_),
    .B1(_04374_),
    .C1(_04372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04377_));
 sky130_fd_sc_hd__a21o_2 _13467_ (.A1(_04372_),
    .A2(_04374_),
    .B1(_04266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04378_));
 sky130_fd_sc_hd__a32oi_2 _13468_ (.A1(_04258_),
    .A2(_04304_),
    .A3(_04305_),
    .B1(_04309_),
    .B2(_04214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04379_));
 sky130_fd_sc_hd__a32o_2 _13469_ (.A1(_04258_),
    .A2(_04304_),
    .A3(_04305_),
    .B1(_04309_),
    .B2(_04214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04380_));
 sky130_fd_sc_hd__nand3_2 _13470_ (.A(_04377_),
    .B(_04378_),
    .C(_04380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04381_));
 sky130_fd_sc_hd__nand3_2 _13471_ (.A(_04375_),
    .B(_04376_),
    .C(_04379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_2 _13472_ (.A(_04381_),
    .B(_04382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04383_));
 sky130_fd_sc_hd__nand3_2 _13473_ (.A(_04314_),
    .B(_04317_),
    .C(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04384_));
 sky130_fd_sc_hd__a21o_2 _13474_ (.A1(_04314_),
    .A2(_04317_),
    .B1(_04383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04385_));
 sky130_fd_sc_hd__and2_2 _13475_ (.A(_04384_),
    .B(_04385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04386_));
 sky130_fd_sc_hd__nand2_2 _13476_ (.A(_04318_),
    .B(_04384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04387_));
 sky130_fd_sc_hd__o211a_2 _13477_ (.A1(_04318_),
    .A2(_04386_),
    .B1(_04387_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00314_));
 sky130_fd_sc_hd__nand3_2 _13478_ (.A(_04316_),
    .B(_04381_),
    .C(_04313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04388_));
 sky130_fd_sc_hd__and4_2 _13479_ (.A(_04381_),
    .B(_04312_),
    .C(_04252_),
    .D(_04251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04389_));
 sky130_fd_sc_hd__a41o_2 _13480_ (.A1(_04327_),
    .A2(_04259_),
    .A3(\a_h[1] ),
    .A4(\a_h[0] ),
    .B1(_04328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04390_));
 sky130_fd_sc_hd__inv_2 _13481_ (.A(_04390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04391_));
 sky130_fd_sc_hd__nand2_2 _13482_ (.A(\a_h[0] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04392_));
 sky130_fd_sc_hd__a21o_2 _13483_ (.A1(_04329_),
    .A2(_04330_),
    .B1(_04392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04393_));
 sky130_fd_sc_hd__a22o_2 _13484_ (.A1(\a_h[0] ),
    .A2(\b_l[9] ),
    .B1(_04327_),
    .B2(_04261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04394_));
 sky130_fd_sc_hd__o21a_2 _13485_ (.A1(_04328_),
    .A2(_04394_),
    .B1(_04393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04395_));
 sky130_fd_sc_hd__inv_2 _13486_ (.A(_04395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04396_));
 sky130_fd_sc_hd__a21o_2 _13487_ (.A1(_04333_),
    .A2(_04366_),
    .B1(_04364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04397_));
 sky130_fd_sc_hd__a21oi_2 _13488_ (.A1(_04333_),
    .A2(_04366_),
    .B1(_04364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04398_));
 sky130_fd_sc_hd__o2bb2ai_2 _13489_ (.A1_N(_04345_),
    .A2_N(_04358_),
    .B1(_04357_),
    .B2(_04353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04399_));
 sky130_fd_sc_hd__a2bb2oi_2 _13490_ (.A1_N(_04353_),
    .A2_N(_04357_),
    .B1(_04358_),
    .B2(_04345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_2 _13491_ (.A(\b_l[5] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_2 _13492_ (.A(\b_l[4] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04402_));
 sky130_fd_sc_hd__nand2_2 _13493_ (.A(\b_l[3] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04403_));
 sky130_fd_sc_hd__nand4_2 _13494_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04404_));
 sky130_fd_sc_hd__a22oi_2 _13495_ (.A1(\b_l[4] ),
    .A2(\a_h[5] ),
    .B1(\a_h[6] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04405_));
 sky130_fd_sc_hd__nand2_2 _13496_ (.A(_04337_),
    .B(_04403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04406_));
 sky130_fd_sc_hd__a22oi_2 _13497_ (.A1(\b_l[5] ),
    .A2(\a_h[4] ),
    .B1(_04404_),
    .B2(_04406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04407_));
 sky130_fd_sc_hd__and3_2 _13498_ (.A(_04404_),
    .B(\a_h[4] ),
    .C(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04408_));
 sky130_fd_sc_hd__a21oi_2 _13499_ (.A1(_04408_),
    .A2(_04406_),
    .B1(_04407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04409_));
 sky130_fd_sc_hd__o21ai_2 _13500_ (.A1(_04348_),
    .A2(_04350_),
    .B1(_04352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04410_));
 sky130_fd_sc_hd__o22a_2 _13501_ (.A1(_02082_),
    .A2(_04134_),
    .B1(_04348_),
    .B2(_04350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04411_));
 sky130_fd_sc_hd__nand2_2 _13502_ (.A(\b_l[1] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_2 _13503_ (.A(\b_l[0] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04413_));
 sky130_fd_sc_hd__a22oi_2 _13504_ (.A1(\b_l[1] ),
    .A2(\a_h[8] ),
    .B1(\a_h[9] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04414_));
 sky130_fd_sc_hd__a22o_2 _13505_ (.A1(\b_l[1] ),
    .A2(\a_h[8] ),
    .B1(\a_h[9] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04415_));
 sky130_fd_sc_hd__nand2_2 _13506_ (.A(\b_l[1] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04416_));
 sky130_fd_sc_hd__nand4_2 _13507_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04417_));
 sky130_fd_sc_hd__o2bb2ai_2 _13508_ (.A1_N(_04412_),
    .A2_N(_04413_),
    .B1(_04416_),
    .B2(_04349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04418_));
 sky130_fd_sc_hd__nor2_2 _13509_ (.A(_09155_),
    .B(_09449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04419_));
 sky130_fd_sc_hd__nand2_2 _13510_ (.A(\b_l[2] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04420_));
 sky130_fd_sc_hd__o221ai_2 _13511_ (.A1(_09155_),
    .A2(_09449_),
    .B1(_04349_),
    .B2(_04416_),
    .C1(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_2 _13512_ (.A(_04418_),
    .B(_04419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04422_));
 sky130_fd_sc_hd__o2111ai_2 _13513_ (.A1(_04349_),
    .A2(_04416_),
    .B1(\b_l[2] ),
    .C1(\a_h[7] ),
    .D1(_04415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04423_));
 sky130_fd_sc_hd__a21oi_2 _13514_ (.A1(_04415_),
    .A2(_04417_),
    .B1(_04419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04424_));
 sky130_fd_sc_hd__o21ai_2 _13515_ (.A1(_09155_),
    .A2(_09449_),
    .B1(_04418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_2 _13516_ (.A1(_04418_),
    .A2(_04420_),
    .B1(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04426_));
 sky130_fd_sc_hd__nand3_2 _13517_ (.A(_04423_),
    .B(_04425_),
    .C(_04410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04427_));
 sky130_fd_sc_hd__nand3_2 _13518_ (.A(_04411_),
    .B(_04421_),
    .C(_04422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04428_));
 sky130_fd_sc_hd__o21ai_2 _13519_ (.A1(_04424_),
    .A2(_04426_),
    .B1(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04429_));
 sky130_fd_sc_hd__o211ai_2 _13520_ (.A1(_04424_),
    .A2(_04426_),
    .B1(_04428_),
    .C1(_04409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04430_));
 sky130_fd_sc_hd__a21o_2 _13521_ (.A1(_04427_),
    .A2(_04428_),
    .B1(_04409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04431_));
 sky130_fd_sc_hd__nand2_2 _13522_ (.A(_04429_),
    .B(_04409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04432_));
 sky130_fd_sc_hd__nand3b_2 _13523_ (.A_N(_04409_),
    .B(_04427_),
    .C(_04428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04433_));
 sky130_fd_sc_hd__nand3_2 _13524_ (.A(_04431_),
    .B(_04399_),
    .C(_04430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04434_));
 sky130_fd_sc_hd__a21oi_2 _13525_ (.A1(_04430_),
    .A2(_04431_),
    .B1(_04399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04435_));
 sky130_fd_sc_hd__nand3_2 _13526_ (.A(_04400_),
    .B(_04432_),
    .C(_04433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04436_));
 sky130_fd_sc_hd__nand2_2 _13527_ (.A(_04434_),
    .B(_04436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04437_));
 sky130_fd_sc_hd__o21ai_2 _13528_ (.A1(_01860_),
    .A2(_04260_),
    .B1(_04324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04438_));
 sky130_fd_sc_hd__nand2_2 _13529_ (.A(\b_l[8] ),
    .B(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_2 _13530_ (.A(\b_l[7] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04440_));
 sky130_fd_sc_hd__nand2_2 _13531_ (.A(\b_l[6] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04441_));
 sky130_fd_sc_hd__nand4_2 _13532_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_2 _13533_ (.A(_04440_),
    .B(_04441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04443_));
 sky130_fd_sc_hd__nand3_2 _13534_ (.A(_04441_),
    .B(\a_h[2] ),
    .C(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04444_));
 sky130_fd_sc_hd__nand3_2 _13535_ (.A(_04440_),
    .B(\a_h[3] ),
    .C(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04445_));
 sky130_fd_sc_hd__nand4_2 _13536_ (.A(_04443_),
    .B(\a_h[1] ),
    .C(\b_l[8] ),
    .D(_04442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04446_));
 sky130_fd_sc_hd__nand3_2 _13537_ (.A(_04439_),
    .B(_04444_),
    .C(_04445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04447_));
 sky130_fd_sc_hd__o21a_2 _13538_ (.A1(_09220_),
    .A2(_09406_),
    .B1(_04338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04448_));
 sky130_fd_sc_hd__o21ai_2 _13539_ (.A1(_09220_),
    .A2(_09406_),
    .B1(_04338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04449_));
 sky130_fd_sc_hd__o2bb2ai_2 _13540_ (.A1_N(_04446_),
    .A2_N(_04447_),
    .B1(_04448_),
    .B2(_04341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04450_));
 sky130_fd_sc_hd__nand4_2 _13541_ (.A(_04342_),
    .B(_04446_),
    .C(_04447_),
    .D(_04449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04451_));
 sky130_fd_sc_hd__a21o_2 _13542_ (.A1(_04450_),
    .A2(_04451_),
    .B1(_04438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04452_));
 sky130_fd_sc_hd__nand3_2 _13543_ (.A(_04438_),
    .B(_04450_),
    .C(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04453_));
 sky130_fd_sc_hd__a22oi_2 _13544_ (.A1(_04321_),
    .A2(_04324_),
    .B1(_04450_),
    .B2(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04454_));
 sky130_fd_sc_hd__and4_2 _13545_ (.A(_04321_),
    .B(_04324_),
    .C(_04450_),
    .D(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04455_));
 sky130_fd_sc_hd__nand2_2 _13546_ (.A(_04452_),
    .B(_04453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04456_));
 sky130_fd_sc_hd__nand3_2 _13547_ (.A(_04434_),
    .B(_04436_),
    .C(_04456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04457_));
 sky130_fd_sc_hd__o2bb2ai_2 _13548_ (.A1_N(_04434_),
    .A2_N(_04436_),
    .B1(_04454_),
    .B2(_04455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04458_));
 sky130_fd_sc_hd__nand2_2 _13549_ (.A(_04437_),
    .B(_04456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04459_));
 sky130_fd_sc_hd__nand3b_2 _13550_ (.A_N(_04456_),
    .B(_04436_),
    .C(_04434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04460_));
 sky130_fd_sc_hd__nand3_2 _13551_ (.A(_04398_),
    .B(_04457_),
    .C(_04458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04461_));
 sky130_fd_sc_hd__a21oi_2 _13552_ (.A1(_04457_),
    .A2(_04458_),
    .B1(_04398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04462_));
 sky130_fd_sc_hd__nand3_2 _13553_ (.A(_04397_),
    .B(_04459_),
    .C(_04460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_2 _13554_ (.A(_04461_),
    .B(_04463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04464_));
 sky130_fd_sc_hd__a21o_2 _13555_ (.A1(_04461_),
    .A2(_04463_),
    .B1(_04395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04465_));
 sky130_fd_sc_hd__and3_2 _13556_ (.A(_04463_),
    .B(_04395_),
    .C(_04461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04466_));
 sky130_fd_sc_hd__nand3_2 _13557_ (.A(_04463_),
    .B(_04395_),
    .C(_04461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04467_));
 sky130_fd_sc_hd__a21o_2 _13558_ (.A1(_04461_),
    .A2(_04463_),
    .B1(_04396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04468_));
 sky130_fd_sc_hd__nand3_2 _13559_ (.A(_04396_),
    .B(_04461_),
    .C(_04463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04469_));
 sky130_fd_sc_hd__a31oi_2 _13560_ (.A1(_04371_),
    .A2(_04319_),
    .A3(_04370_),
    .B1(_04265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04470_));
 sky130_fd_sc_hd__a32oi_2 _13561_ (.A1(_04320_),
    .A2(_04368_),
    .A3(_04369_),
    .B1(_04372_),
    .B2(_04266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04471_));
 sky130_fd_sc_hd__o211ai_2 _13562_ (.A1(_04373_),
    .A2(_04470_),
    .B1(_04469_),
    .C1(_04468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04472_));
 sky130_fd_sc_hd__a211o_2 _13563_ (.A1(_04396_),
    .A2(_04464_),
    .B1(_04470_),
    .C1(_04373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04473_));
 sky130_fd_sc_hd__nand3_2 _13564_ (.A(_04465_),
    .B(_04467_),
    .C(_04471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04474_));
 sky130_fd_sc_hd__inv_2 _13565_ (.A(_04474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04475_));
 sky130_fd_sc_hd__nand2_2 _13566_ (.A(_04472_),
    .B(_04474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04476_));
 sky130_fd_sc_hd__nand2_2 _13567_ (.A(_04382_),
    .B(_04476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04477_));
 sky130_fd_sc_hd__nand3b_2 _13568_ (.A_N(_04382_),
    .B(_04472_),
    .C(_04474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04478_));
 sky130_fd_sc_hd__a21oi_2 _13569_ (.A1(_04477_),
    .A2(_04478_),
    .B1(_04389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04479_));
 sky130_fd_sc_hd__a21o_2 _13570_ (.A1(_04389_),
    .A2(_04477_),
    .B1(_04479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04480_));
 sky130_fd_sc_hd__nand3_2 _13571_ (.A(_04387_),
    .B(_04388_),
    .C(_04480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04481_));
 sky130_fd_sc_hd__a221o_2 _13572_ (.A1(_04389_),
    .A2(_04477_),
    .B1(_04387_),
    .B2(_04388_),
    .C1(_04479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04482_));
 sky130_fd_sc_hd__and3_2 _13573_ (.A(_09690_),
    .B(_04481_),
    .C(_04482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00315_));
 sky130_fd_sc_hd__a21oi_2 _13574_ (.A1(_04314_),
    .A2(_04476_),
    .B1(_04388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04483_));
 sky130_fd_sc_hd__a21oi_2 _13575_ (.A1(_04389_),
    .A2(_04477_),
    .B1(_04483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04484_));
 sky130_fd_sc_hd__o21ai_2 _13576_ (.A1(_04387_),
    .A2(_04479_),
    .B1(_04484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04485_));
 sky130_fd_sc_hd__a32oi_2 _13577_ (.A1(_04431_),
    .A2(_04399_),
    .A3(_04430_),
    .B1(_04452_),
    .B2(_04453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04486_));
 sky130_fd_sc_hd__a21oi_2 _13578_ (.A1(_04434_),
    .A2(_04456_),
    .B1(_04435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04487_));
 sky130_fd_sc_hd__o21ai_2 _13579_ (.A1(_01871_),
    .A2(_04260_),
    .B1(_04446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_2 _13580_ (.A(\b_l[7] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04489_));
 sky130_fd_sc_hd__nand2_2 _13581_ (.A(\b_l[6] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_2 _13582_ (.A(_04489_),
    .B(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04491_));
 sky130_fd_sc_hd__o2111ai_2 _13583_ (.A1(_01888_),
    .A2(_04260_),
    .B1(\b_l[8] ),
    .C1(\a_h[2] ),
    .D1(_04491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04492_));
 sky130_fd_sc_hd__nand3_2 _13584_ (.A(_04490_),
    .B(\a_h[3] ),
    .C(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04493_));
 sky130_fd_sc_hd__nand3_2 _13585_ (.A(_04489_),
    .B(\a_h[4] ),
    .C(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04494_));
 sky130_fd_sc_hd__o211ai_2 _13586_ (.A1(_09264_),
    .A2(_09395_),
    .B1(_04493_),
    .C1(_04494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04495_));
 sky130_fd_sc_hd__o22a_2 _13587_ (.A1(_09220_),
    .A2(_09417_),
    .B1(_04337_),
    .B2(_04403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04496_));
 sky130_fd_sc_hd__a21oi_2 _13588_ (.A1(_04401_),
    .A2(_04404_),
    .B1(_04405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04497_));
 sky130_fd_sc_hd__o2bb2ai_2 _13589_ (.A1_N(_04492_),
    .A2_N(_04495_),
    .B1(_04496_),
    .B2(_04405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04498_));
 sky130_fd_sc_hd__nand3_2 _13590_ (.A(_04492_),
    .B(_04495_),
    .C(_04497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04499_));
 sky130_fd_sc_hd__inv_2 _13591_ (.A(_04499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04500_));
 sky130_fd_sc_hd__nand2_2 _13592_ (.A(_04488_),
    .B(_04498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04501_));
 sky130_fd_sc_hd__a21o_2 _13593_ (.A1(_04498_),
    .A2(_04499_),
    .B1(_04488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04502_));
 sky130_fd_sc_hd__o21ai_2 _13594_ (.A1(_04500_),
    .A2(_04501_),
    .B1(_04502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04503_));
 sky130_fd_sc_hd__o2bb2ai_2 _13595_ (.A1_N(_04409_),
    .A2_N(_04428_),
    .B1(_04426_),
    .B2(_04424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04504_));
 sky130_fd_sc_hd__a21boi_2 _13596_ (.A1(_04409_),
    .A2(_04428_),
    .B1_N(_04427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04505_));
 sky130_fd_sc_hd__nand2_2 _13597_ (.A(\b_l[5] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04506_));
 sky130_fd_sc_hd__nand2_2 _13598_ (.A(\b_l[3] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04507_));
 sky130_fd_sc_hd__nand4_2 _13599_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[6] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04508_));
 sky130_fd_sc_hd__a22oi_2 _13600_ (.A1(\b_l[4] ),
    .A2(\a_h[6] ),
    .B1(\a_h[7] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_2 _13601_ (.A(_04402_),
    .B(_04507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04510_));
 sky130_fd_sc_hd__o2bb2a_2 _13602_ (.A1_N(_04508_),
    .A2_N(_04510_),
    .B1(_09220_),
    .B2(_09428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04511_));
 sky130_fd_sc_hd__and4_2 _13603_ (.A(_04510_),
    .B(\a_h[5] ),
    .C(\b_l[5] ),
    .D(_04508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04512_));
 sky130_fd_sc_hd__a21o_2 _13604_ (.A1(_04508_),
    .A2(_04510_),
    .B1(_04506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04513_));
 sky130_fd_sc_hd__o21ai_2 _13605_ (.A1(_04402_),
    .A2(_04507_),
    .B1(_04506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04514_));
 sky130_fd_sc_hd__o211ai_2 _13606_ (.A1(_09220_),
    .A2(_09428_),
    .B1(_04508_),
    .C1(_04510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04515_));
 sky130_fd_sc_hd__o21ai_2 _13607_ (.A1(_04509_),
    .A2(_04514_),
    .B1(_04513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04516_));
 sky130_fd_sc_hd__and2_2 _13608_ (.A(\b_l[2] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04517_));
 sky130_fd_sc_hd__nand2_2 _13609_ (.A(\b_l[2] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_2 _13610_ (.A(\b_l[0] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04519_));
 sky130_fd_sc_hd__a22oi_2 _13611_ (.A1(\b_l[1] ),
    .A2(\a_h[9] ),
    .B1(\a_h[10] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_2 _13612_ (.A(_04416_),
    .B(_04519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04521_));
 sky130_fd_sc_hd__nand4_2 _13613_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04522_));
 sky130_fd_sc_hd__nand2_2 _13614_ (.A(_04521_),
    .B(_04522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04523_));
 sky130_fd_sc_hd__a21o_2 _13615_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04524_));
 sky130_fd_sc_hd__nand4_2 _13616_ (.A(_04521_),
    .B(_04522_),
    .C(\b_l[2] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04525_));
 sky130_fd_sc_hd__nand2_2 _13617_ (.A(_04417_),
    .B(_04420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04526_));
 sky130_fd_sc_hd__o21ai_2 _13618_ (.A1(_04420_),
    .A2(_04414_),
    .B1(_04417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04527_));
 sky130_fd_sc_hd__o22a_2 _13619_ (.A1(_04349_),
    .A2(_04416_),
    .B1(_04420_),
    .B2(_04414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04528_));
 sky130_fd_sc_hd__and3_2 _13620_ (.A(_04524_),
    .B(_04525_),
    .C(_04527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04529_));
 sky130_fd_sc_hd__nand3_2 _13621_ (.A(_04524_),
    .B(_04525_),
    .C(_04527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04530_));
 sky130_fd_sc_hd__o211ai_2 _13622_ (.A1(_09155_),
    .A2(_09460_),
    .B1(_04521_),
    .C1(_04522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04531_));
 sky130_fd_sc_hd__a21o_2 _13623_ (.A1(_04521_),
    .A2(_04522_),
    .B1(_04518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04532_));
 sky130_fd_sc_hd__a22oi_2 _13624_ (.A1(_04415_),
    .A2(_04526_),
    .B1(_04523_),
    .B2(_04517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04533_));
 sky130_fd_sc_hd__nand3_2 _13625_ (.A(_04528_),
    .B(_04531_),
    .C(_04532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_2 _13626_ (.A(_04530_),
    .B(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04535_));
 sky130_fd_sc_hd__o211a_2 _13627_ (.A1(_04511_),
    .A2(_04512_),
    .B1(_04530_),
    .C1(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04536_));
 sky130_fd_sc_hd__o2111ai_2 _13628_ (.A1(_04514_),
    .A2(_04509_),
    .B1(_04513_),
    .C1(_04530_),
    .D1(_04534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_2 _13629_ (.A(_04535_),
    .B(_04516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04538_));
 sky130_fd_sc_hd__o21ai_2 _13630_ (.A1(_04511_),
    .A2(_04512_),
    .B1(_04535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04539_));
 sky130_fd_sc_hd__a22oi_2 _13631_ (.A1(_04513_),
    .A2(_04515_),
    .B1(_04533_),
    .B2(_04531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_2 _13632_ (.A(_04540_),
    .B(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04541_));
 sky130_fd_sc_hd__nand2_2 _13633_ (.A(_04505_),
    .B(_04538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04542_));
 sky130_fd_sc_hd__nand3_2 _13634_ (.A(_04505_),
    .B(_04537_),
    .C(_04538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04543_));
 sky130_fd_sc_hd__nand3_2 _13635_ (.A(_04539_),
    .B(_04541_),
    .C(_04504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_2 _13636_ (.A(_04543_),
    .B(_04544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04545_));
 sky130_fd_sc_hd__o211ai_2 _13637_ (.A1(_04536_),
    .A2(_04542_),
    .B1(_04544_),
    .C1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04546_));
 sky130_fd_sc_hd__a21o_2 _13638_ (.A1(_04543_),
    .A2(_04544_),
    .B1(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04547_));
 sky130_fd_sc_hd__o2111ai_2 _13639_ (.A1(_04500_),
    .A2(_04501_),
    .B1(_04502_),
    .C1(_04543_),
    .D1(_04544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04548_));
 sky130_fd_sc_hd__nand2_2 _13640_ (.A(_04503_),
    .B(_04545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_2 _13641_ (.A(_04546_),
    .B(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04550_));
 sky130_fd_sc_hd__o211ai_2 _13642_ (.A1(_04435_),
    .A2(_04486_),
    .B1(_04546_),
    .C1(_04547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04551_));
 sky130_fd_sc_hd__and3_2 _13643_ (.A(_04549_),
    .B(_04487_),
    .C(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04552_));
 sky130_fd_sc_hd__nand3_2 _13644_ (.A(_04549_),
    .B(_04487_),
    .C(_04548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04553_));
 sky130_fd_sc_hd__and2_2 _13645_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04554_));
 sky130_fd_sc_hd__nand2_2 _13646_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04555_));
 sky130_fd_sc_hd__and3_2 _13647_ (.A(\a_h[0] ),
    .B(\a_h[1] ),
    .C(_04554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04556_));
 sky130_fd_sc_hd__a22oi_2 _13648_ (.A1(\a_h[0] ),
    .A2(\b_l[10] ),
    .B1(\a_h[1] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04557_));
 sky130_fd_sc_hd__a31o_2 _13649_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04554_),
    .B1(_04557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04558_));
 sky130_fd_sc_hd__a21bo_2 _13650_ (.A1(_04438_),
    .A2(_04450_),
    .B1_N(_04451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04559_));
 sky130_fd_sc_hd__inv_2 _13651_ (.A(_04559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04560_));
 sky130_fd_sc_hd__o21a_2 _13652_ (.A1(_04556_),
    .A2(_04557_),
    .B1(_04560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04561_));
 sky130_fd_sc_hd__nor2_2 _13653_ (.A(_04558_),
    .B(_04560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04562_));
 sky130_fd_sc_hd__a311o_2 _13654_ (.A1(\a_h[0] ),
    .A2(\a_h[1] ),
    .A3(_04554_),
    .B1(_04557_),
    .C1(_04560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_2 _13655_ (.A(_04558_),
    .B(_04559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04564_));
 sky130_fd_sc_hd__inv_2 _13656_ (.A(_04564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04565_));
 sky130_fd_sc_hd__o2bb2ai_2 _13657_ (.A1_N(_04551_),
    .A2_N(_04553_),
    .B1(_04561_),
    .B2(_04562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04566_));
 sky130_fd_sc_hd__nand2_2 _13658_ (.A(_04551_),
    .B(_04564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04567_));
 sky130_fd_sc_hd__nand3_2 _13659_ (.A(_04551_),
    .B(_04553_),
    .C(_04564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04568_));
 sky130_fd_sc_hd__a21o_2 _13660_ (.A1(_04395_),
    .A2(_04461_),
    .B1(_04462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04569_));
 sky130_fd_sc_hd__a21oi_2 _13661_ (.A1(_04566_),
    .A2(_04568_),
    .B1(_04569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04570_));
 sky130_fd_sc_hd__a21o_2 _13662_ (.A1(_04566_),
    .A2(_04568_),
    .B1(_04569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04571_));
 sky130_fd_sc_hd__o211a_2 _13663_ (.A1(_04552_),
    .A2(_04567_),
    .B1(_04566_),
    .C1(_04569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04572_));
 sky130_fd_sc_hd__o211ai_2 _13664_ (.A1(_04552_),
    .A2(_04567_),
    .B1(_04566_),
    .C1(_04569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04573_));
 sky130_fd_sc_hd__o22ai_2 _13665_ (.A1(_04391_),
    .A2(_04392_),
    .B1(_04570_),
    .B2(_04572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04574_));
 sky130_fd_sc_hd__nand3b_2 _13666_ (.A_N(_04393_),
    .B(_04571_),
    .C(_04573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04575_));
 sky130_fd_sc_hd__o211ai_2 _13667_ (.A1(_04391_),
    .A2(_04392_),
    .B1(_04571_),
    .C1(_04573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04576_));
 sky130_fd_sc_hd__o21bai_2 _13668_ (.A1(_04570_),
    .A2(_04572_),
    .B1_N(_04393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04577_));
 sky130_fd_sc_hd__o211ai_2 _13669_ (.A1(_04466_),
    .A2(_04473_),
    .B1(_04576_),
    .C1(_04577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04578_));
 sky130_fd_sc_hd__nand3_2 _13670_ (.A(_04574_),
    .B(_04575_),
    .C(_04475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04579_));
 sky130_fd_sc_hd__o2bb2ai_2 _13671_ (.A1_N(_04578_),
    .A2_N(_04579_),
    .B1(_04382_),
    .B2(_04476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04580_));
 sky130_fd_sc_hd__a21o_2 _13672_ (.A1(_04576_),
    .A2(_04577_),
    .B1(_04478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04581_));
 sky130_fd_sc_hd__a21o_2 _13673_ (.A1(_04580_),
    .A2(_04581_),
    .B1(_04485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04582_));
 sky130_fd_sc_hd__nand2_2 _13674_ (.A(_04485_),
    .B(_04580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04583_));
 sky130_fd_sc_hd__and3_2 _13675_ (.A(_09690_),
    .B(_04582_),
    .C(_04583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00316_));
 sky130_fd_sc_hd__nand2_2 _13676_ (.A(_04553_),
    .B(_04565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04584_));
 sky130_fd_sc_hd__o21ai_2 _13677_ (.A1(_04487_),
    .A2(_04550_),
    .B1(_04584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04585_));
 sky130_fd_sc_hd__a32oi_2 _13678_ (.A1(_04505_),
    .A2(_04537_),
    .A3(_04538_),
    .B1(_04544_),
    .B2(_04503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04586_));
 sky130_fd_sc_hd__o2bb2ai_2 _13679_ (.A1_N(_04503_),
    .A2_N(_04544_),
    .B1(_04542_),
    .B2(_04536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04587_));
 sky130_fd_sc_hd__a21boi_2 _13680_ (.A1(_04534_),
    .A2(_04516_),
    .B1_N(_04530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04588_));
 sky130_fd_sc_hd__o2bb2a_2 _13681_ (.A1_N(\b_l[2] ),
    .A2_N(\a_h[8] ),
    .B1(_04416_),
    .B2(_04519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04589_));
 sky130_fd_sc_hd__o21ai_2 _13682_ (.A1(_04518_),
    .A2(_04520_),
    .B1(_04522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04590_));
 sky130_fd_sc_hd__and2_2 _13683_ (.A(\b_l[2] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_2 _13684_ (.A(\b_l[2] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2_2 _13685_ (.A(\b_l[1] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_2 _13686_ (.A(\b_l[0] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04594_));
 sky130_fd_sc_hd__a22oi_2 _13687_ (.A1(\b_l[1] ),
    .A2(\a_h[10] ),
    .B1(\a_h[11] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_2 _13688_ (.A(_04593_),
    .B(_04594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04596_));
 sky130_fd_sc_hd__nand4_2 _13689_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04597_));
 sky130_fd_sc_hd__o21ai_2 _13690_ (.A1(_02362_),
    .A2(_04134_),
    .B1(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04598_));
 sky130_fd_sc_hd__o221a_2 _13691_ (.A1(_09155_),
    .A2(_09471_),
    .B1(_02362_),
    .B2(_04134_),
    .C1(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04599_));
 sky130_fd_sc_hd__o221ai_2 _13692_ (.A1(_09155_),
    .A2(_09471_),
    .B1(_02362_),
    .B2(_04134_),
    .C1(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04600_));
 sky130_fd_sc_hd__a21o_2 _13693_ (.A1(_04596_),
    .A2(_04597_),
    .B1(_04592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04601_));
 sky130_fd_sc_hd__o2111ai_2 _13694_ (.A1(_02362_),
    .A2(_04134_),
    .B1(\b_l[2] ),
    .C1(\a_h[9] ),
    .D1(_04596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04602_));
 sky130_fd_sc_hd__a21o_2 _13695_ (.A1(_04596_),
    .A2(_04597_),
    .B1(_04591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04603_));
 sky130_fd_sc_hd__nand3_2 _13696_ (.A(_04603_),
    .B(_04590_),
    .C(_04602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04604_));
 sky130_fd_sc_hd__o2bb2ai_2 _13697_ (.A1_N(_04591_),
    .A2_N(_04598_),
    .B1(_04520_),
    .B2(_04589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04605_));
 sky130_fd_sc_hd__o211ai_2 _13698_ (.A1(_04520_),
    .A2(_04589_),
    .B1(_04600_),
    .C1(_04601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_2 _13699_ (.A(\b_l[5] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04607_));
 sky130_fd_sc_hd__a22oi_2 _13700_ (.A1(\b_l[4] ),
    .A2(\a_h[7] ),
    .B1(\a_h[8] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_2 _13701_ (.A(_02082_),
    .B(_04182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04609_));
 sky130_fd_sc_hd__nand4_2 _13702_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04610_));
 sky130_fd_sc_hd__o211a_2 _13703_ (.A1(_04608_),
    .A2(_04609_),
    .B1(\b_l[5] ),
    .C1(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04611_));
 sky130_fd_sc_hd__a211oi_2 _13704_ (.A1(\b_l[5] ),
    .A2(\a_h[6] ),
    .B1(_04608_),
    .C1(_04609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04612_));
 sky130_fd_sc_hd__a41o_2 _13705_ (.A1(\b_l[3] ),
    .A2(\b_l[4] ),
    .A3(\a_h[7] ),
    .A4(\a_h[8] ),
    .B1(_04607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04613_));
 sky130_fd_sc_hd__and4b_2 _13706_ (.A_N(_04608_),
    .B(_04610_),
    .C(\b_l[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04614_));
 sky130_fd_sc_hd__o22a_2 _13707_ (.A1(_09220_),
    .A2(_09439_),
    .B1(_04608_),
    .B2(_04609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04615_));
 sky130_fd_sc_hd__o21ai_2 _13708_ (.A1(_04608_),
    .A2(_04609_),
    .B1(_04607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04616_));
 sky130_fd_sc_hd__o21ai_2 _13709_ (.A1(_04608_),
    .A2(_04613_),
    .B1(_04616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04617_));
 sky130_fd_sc_hd__o21a_2 _13710_ (.A1(_04608_),
    .A2(_04613_),
    .B1(_04616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04618_));
 sky130_fd_sc_hd__o221a_2 _13711_ (.A1(_04599_),
    .A2(_04605_),
    .B1(_04614_),
    .B2(_04615_),
    .C1(_04604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04619_));
 sky130_fd_sc_hd__nand3_2 _13712_ (.A(_04604_),
    .B(_04606_),
    .C(_04617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04620_));
 sky130_fd_sc_hd__o2bb2ai_2 _13713_ (.A1_N(_04604_),
    .A2_N(_04606_),
    .B1(_04611_),
    .B2(_04612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04621_));
 sky130_fd_sc_hd__o211ai_2 _13714_ (.A1(_04599_),
    .A2(_04605_),
    .B1(_04618_),
    .C1(_04604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04622_));
 sky130_fd_sc_hd__o2bb2ai_2 _13715_ (.A1_N(_04604_),
    .A2_N(_04606_),
    .B1(_04614_),
    .B2(_04615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04623_));
 sky130_fd_sc_hd__nand2_2 _13716_ (.A(_04621_),
    .B(_04588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04624_));
 sky130_fd_sc_hd__nand3_2 _13717_ (.A(_04621_),
    .B(_04588_),
    .C(_04620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04625_));
 sky130_fd_sc_hd__o211ai_2 _13718_ (.A1(_04529_),
    .A2(_04540_),
    .B1(_04622_),
    .C1(_04623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04626_));
 sky130_fd_sc_hd__o31a_2 _13719_ (.A1(_09406_),
    .A2(_09417_),
    .A3(_04260_),
    .B1(_04492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04627_));
 sky130_fd_sc_hd__o21ai_2 _13720_ (.A1(_01888_),
    .A2(_04260_),
    .B1(_04492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04628_));
 sky130_fd_sc_hd__a21o_2 _13721_ (.A1(_04506_),
    .A2(_04508_),
    .B1(_04509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04629_));
 sky130_fd_sc_hd__a21oi_2 _13722_ (.A1(_04506_),
    .A2(_04508_),
    .B1(_04509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_2 _13723_ (.A(\b_l[8] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04631_));
 sky130_fd_sc_hd__nand2_2 _13724_ (.A(\b_l[6] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04632_));
 sky130_fd_sc_hd__a22oi_2 _13725_ (.A1(\b_l[7] ),
    .A2(\a_h[4] ),
    .B1(\a_h[5] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04633_));
 sky130_fd_sc_hd__a22o_2 _13726_ (.A1(\b_l[7] ),
    .A2(\a_h[4] ),
    .B1(\a_h[5] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_2 _13727_ (.A(\b_l[7] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04635_));
 sky130_fd_sc_hd__and4_2 _13728_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04636_));
 sky130_fd_sc_hd__a41o_2 _13729_ (.A1(\b_l[6] ),
    .A2(\b_l[7] ),
    .A3(\a_h[4] ),
    .A4(\a_h[5] ),
    .B1(_04631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04637_));
 sky130_fd_sc_hd__o21ai_2 _13730_ (.A1(_04633_),
    .A2(_04636_),
    .B1(_04631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04638_));
 sky130_fd_sc_hd__o21bai_2 _13731_ (.A1(_04633_),
    .A2(_04636_),
    .B1_N(_04631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04639_));
 sky130_fd_sc_hd__o221ai_2 _13732_ (.A1(_09264_),
    .A2(_09406_),
    .B1(_04490_),
    .B2(_04635_),
    .C1(_04634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04640_));
 sky130_fd_sc_hd__o211ai_2 _13733_ (.A1(_04637_),
    .A2(_04633_),
    .B1(_04630_),
    .C1(_04638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04641_));
 sky130_fd_sc_hd__nand3_2 _13734_ (.A(_04639_),
    .B(_04640_),
    .C(_04629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04642_));
 sky130_fd_sc_hd__a21oi_2 _13735_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04643_));
 sky130_fd_sc_hd__a21o_2 _13736_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04644_));
 sky130_fd_sc_hd__and3_2 _13737_ (.A(_04628_),
    .B(_04641_),
    .C(_04642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04645_));
 sky130_fd_sc_hd__nand3_2 _13738_ (.A(_04628_),
    .B(_04641_),
    .C(_04642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04646_));
 sky130_fd_sc_hd__a21oi_2 _13739_ (.A1(_04641_),
    .A2(_04642_),
    .B1(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04647_));
 sky130_fd_sc_hd__and3_2 _13740_ (.A(_04627_),
    .B(_04641_),
    .C(_04642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04648_));
 sky130_fd_sc_hd__nand2_2 _13741_ (.A(_04644_),
    .B(_04646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04649_));
 sky130_fd_sc_hd__o211ai_2 _13742_ (.A1(_04619_),
    .A2(_04624_),
    .B1(_04626_),
    .C1(_04649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04650_));
 sky130_fd_sc_hd__o2bb2ai_2 _13743_ (.A1_N(_04625_),
    .A2_N(_04626_),
    .B1(_04647_),
    .B2(_04648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04651_));
 sky130_fd_sc_hd__o2bb2ai_2 _13744_ (.A1_N(_04626_),
    .A2_N(_04649_),
    .B1(_04619_),
    .B2(_04624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04652_));
 sky130_fd_sc_hd__a21boi_2 _13745_ (.A1(_04626_),
    .A2(_04649_),
    .B1_N(_04625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04653_));
 sky130_fd_sc_hd__and3_2 _13746_ (.A(_04587_),
    .B(_04650_),
    .C(_04651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04654_));
 sky130_fd_sc_hd__nand3_2 _13747_ (.A(_04587_),
    .B(_04650_),
    .C(_04651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04655_));
 sky130_fd_sc_hd__o211ai_2 _13748_ (.A1(_04647_),
    .A2(_04648_),
    .B1(_04625_),
    .C1(_04626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04656_));
 sky130_fd_sc_hd__inv_2 _13749_ (.A(_04656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04657_));
 sky130_fd_sc_hd__o2bb2ai_2 _13750_ (.A1_N(_04625_),
    .A2_N(_04626_),
    .B1(_04643_),
    .B2(_04645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_2 _13751_ (.A(_04586_),
    .B(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04659_));
 sky130_fd_sc_hd__nand3_2 _13752_ (.A(_04586_),
    .B(_04656_),
    .C(_04658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04660_));
 sky130_fd_sc_hd__nand2_2 _13753_ (.A(\a_h[0] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04661_));
 sky130_fd_sc_hd__a22oi_2 _13754_ (.A1(\b_l[10] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04662_));
 sky130_fd_sc_hd__a22o_2 _13755_ (.A1(\b_l[10] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04663_));
 sky130_fd_sc_hd__nand4_2 _13756_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04664_));
 sky130_fd_sc_hd__o221a_2 _13757_ (.A1(_09177_),
    .A2(_09308_),
    .B1(_01860_),
    .B2(_04555_),
    .C1(_04663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04665_));
 sky130_fd_sc_hd__a21oi_2 _13758_ (.A1(_04663_),
    .A2(_04664_),
    .B1(_04661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04666_));
 sky130_fd_sc_hd__o2111a_2 _13759_ (.A1(_04665_),
    .A2(_04666_),
    .B1(\a_h[0] ),
    .C1(\a_h[1] ),
    .D1(_04554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04667_));
 sky130_fd_sc_hd__o21ai_2 _13760_ (.A1(_04665_),
    .A2(_04666_),
    .B1(_04556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04668_));
 sky130_fd_sc_hd__a31o_2 _13761_ (.A1(_04661_),
    .A2(_04663_),
    .A3(_04664_),
    .B1(_04556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04669_));
 sky130_fd_sc_hd__o21ai_2 _13762_ (.A1(_04666_),
    .A2(_04669_),
    .B1(_04668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04670_));
 sky130_fd_sc_hd__a21o_2 _13763_ (.A1(_04488_),
    .A2(_04498_),
    .B1(_04500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04671_));
 sky130_fd_sc_hd__a21oi_2 _13764_ (.A1(_04488_),
    .A2(_04498_),
    .B1(_04500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04672_));
 sky130_fd_sc_hd__o211a_2 _13765_ (.A1(_04666_),
    .A2(_04669_),
    .B1(_04668_),
    .C1(_04671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04673_));
 sky130_fd_sc_hd__and3_2 _13766_ (.A(_04499_),
    .B(_04501_),
    .C(_04670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04674_));
 sky130_fd_sc_hd__and2_2 _13767_ (.A(_04671_),
    .B(_04670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04675_));
 sky130_fd_sc_hd__o211a_2 _13768_ (.A1(_04669_),
    .A2(_04666_),
    .B1(_04668_),
    .C1(_04672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04676_));
 sky130_fd_sc_hd__xnor2_2 _13769_ (.A(_04670_),
    .B(_04671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04677_));
 sky130_fd_sc_hd__o211ai_2 _13770_ (.A1(_04675_),
    .A2(_04676_),
    .B1(_04655_),
    .C1(_04660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04678_));
 sky130_fd_sc_hd__o2bb2ai_2 _13771_ (.A1_N(_04655_),
    .A2_N(_04660_),
    .B1(_04673_),
    .B2(_04674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04679_));
 sky130_fd_sc_hd__o2111a_2 _13772_ (.A1(_04487_),
    .A2(_04550_),
    .B1(_04584_),
    .C1(_04678_),
    .D1(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04680_));
 sky130_fd_sc_hd__o2111ai_2 _13773_ (.A1(_04487_),
    .A2(_04550_),
    .B1(_04584_),
    .C1(_04678_),
    .D1(_04679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04681_));
 sky130_fd_sc_hd__a31oi_2 _13774_ (.A1(_04586_),
    .A2(_04656_),
    .A3(_04658_),
    .B1(_04677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04682_));
 sky130_fd_sc_hd__nand2_2 _13775_ (.A(_04682_),
    .B(_04655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04683_));
 sky130_fd_sc_hd__inv_2 _13776_ (.A(_04683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04684_));
 sky130_fd_sc_hd__o2bb2ai_2 _13777_ (.A1_N(_04655_),
    .A2_N(_04660_),
    .B1(_04675_),
    .B2(_04676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2_2 _13778_ (.A(_04585_),
    .B(_04685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04686_));
 sky130_fd_sc_hd__nand3_2 _13779_ (.A(_04585_),
    .B(_04683_),
    .C(_04685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04687_));
 sky130_fd_sc_hd__o2bb2ai_2 _13780_ (.A1_N(_04681_),
    .A2_N(_04687_),
    .B1(_04558_),
    .B2(_04560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04688_));
 sky130_fd_sc_hd__nand3_2 _13781_ (.A(_04687_),
    .B(_04562_),
    .C(_04681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04689_));
 sky130_fd_sc_hd__o21ai_2 _13782_ (.A1(_04393_),
    .A2(_04570_),
    .B1(_04573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04690_));
 sky130_fd_sc_hd__a21oi_2 _13783_ (.A1(_04688_),
    .A2(_04689_),
    .B1(_04690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04691_));
 sky130_fd_sc_hd__a21o_2 _13784_ (.A1(_04688_),
    .A2(_04689_),
    .B1(_04690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04692_));
 sky130_fd_sc_hd__nand3_2 _13785_ (.A(_04690_),
    .B(_04689_),
    .C(_04688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04693_));
 sky130_fd_sc_hd__a32oi_2 _13786_ (.A1(_04475_),
    .A2(_04574_),
    .A3(_04575_),
    .B1(_04692_),
    .B2(_04693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04694_));
 sky130_fd_sc_hd__a21bo_2 _13787_ (.A1(_04692_),
    .A2(_04693_),
    .B1_N(_04579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04695_));
 sky130_fd_sc_hd__a211o_2 _13788_ (.A1(_04576_),
    .A2(_04577_),
    .B1(_04474_),
    .C1(_04691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04696_));
 sky130_fd_sc_hd__a41o_2 _13789_ (.A1(_04475_),
    .A2(_04574_),
    .A3(_04575_),
    .A4(_04692_),
    .B1(_04694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04697_));
 sky130_fd_sc_hd__and3_2 _13790_ (.A(_04581_),
    .B(_04583_),
    .C(_04697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04698_));
 sky130_fd_sc_hd__a21o_2 _13791_ (.A1(_04581_),
    .A2(_04583_),
    .B1(_04694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04699_));
 sky130_fd_sc_hd__nor3b_2 _13792_ (.A(rst),
    .B(_04698_),
    .C_N(_04699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00317_));
 sky130_fd_sc_hd__a31oi_2 _13793_ (.A1(_04585_),
    .A2(_04683_),
    .A3(_04685_),
    .B1(_04563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04700_));
 sky130_fd_sc_hd__o2bb2ai_2 _13794_ (.A1_N(_04563_),
    .A2_N(_04681_),
    .B1(_04684_),
    .B2(_04686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04701_));
 sky130_fd_sc_hd__o2bb2ai_2 _13795_ (.A1_N(_04655_),
    .A2_N(_04677_),
    .B1(_04657_),
    .B2(_04659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04702_));
 sky130_fd_sc_hd__o22a_2 _13796_ (.A1(_09220_),
    .A2(_09439_),
    .B1(_02082_),
    .B2(_04182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04703_));
 sky130_fd_sc_hd__o21ai_2 _13797_ (.A1(_02082_),
    .A2(_04182_),
    .B1(_04607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_2 _13798_ (.A1(_04607_),
    .A2(_04610_),
    .B1(_04608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_2 _13799_ (.A(\b_l[8] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_2 _13800_ (.A(\b_l[7] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04707_));
 sky130_fd_sc_hd__nand2_2 _13801_ (.A(\b_l[6] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04708_));
 sky130_fd_sc_hd__and4_2 _13802_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04709_));
 sky130_fd_sc_hd__nand4_2 _13803_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_2 _13804_ (.A(_04635_),
    .B(_04708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04711_));
 sky130_fd_sc_hd__o221ai_2 _13805_ (.A1(_09264_),
    .A2(_09417_),
    .B1(_04632_),
    .B2(_04707_),
    .C1(_04711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04712_));
 sky130_fd_sc_hd__a21o_2 _13806_ (.A1(_04710_),
    .A2(_04711_),
    .B1(_04706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04713_));
 sky130_fd_sc_hd__o2111ai_2 _13807_ (.A1(_04632_),
    .A2(_04707_),
    .B1(\b_l[8] ),
    .C1(\a_h[4] ),
    .D1(_04711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04714_));
 sky130_fd_sc_hd__nand3_2 _13808_ (.A(_04708_),
    .B(\a_h[5] ),
    .C(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04715_));
 sky130_fd_sc_hd__nand3_2 _13809_ (.A(_04635_),
    .B(\a_h[6] ),
    .C(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04716_));
 sky130_fd_sc_hd__o211ai_2 _13810_ (.A1(_09264_),
    .A2(_09417_),
    .B1(_04715_),
    .C1(_04716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04717_));
 sky130_fd_sc_hd__a21oi_2 _13811_ (.A1(_04714_),
    .A2(_04717_),
    .B1(_04705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04718_));
 sky130_fd_sc_hd__o211ai_2 _13812_ (.A1(_04608_),
    .A2(_04703_),
    .B1(_04712_),
    .C1(_04713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04719_));
 sky130_fd_sc_hd__nand3_2 _13813_ (.A(_04704_),
    .B(_04714_),
    .C(_04717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04720_));
 sky130_fd_sc_hd__nand3_2 _13814_ (.A(_04705_),
    .B(_04714_),
    .C(_04717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04721_));
 sky130_fd_sc_hd__o32a_2 _13815_ (.A1(_09264_),
    .A2(_09406_),
    .A3(_04633_),
    .B1(_04635_),
    .B2(_04490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04722_));
 sky130_fd_sc_hd__a21oi_2 _13816_ (.A1(_04719_),
    .A2(_04721_),
    .B1(_04722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04723_));
 sky130_fd_sc_hd__a21o_2 _13817_ (.A1(_04719_),
    .A2(_04721_),
    .B1(_04722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04724_));
 sky130_fd_sc_hd__nand2_2 _13818_ (.A(_04722_),
    .B(_04721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04725_));
 sky130_fd_sc_hd__and3_2 _13819_ (.A(_04719_),
    .B(_04721_),
    .C(_04722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04726_));
 sky130_fd_sc_hd__o21ai_2 _13820_ (.A1(_04718_),
    .A2(_04725_),
    .B1(_04724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04727_));
 sky130_fd_sc_hd__a2bb2oi_2 _13821_ (.A1_N(_04599_),
    .A2_N(_04605_),
    .B1(_04617_),
    .B2(_04604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04728_));
 sky130_fd_sc_hd__o2bb2ai_2 _13822_ (.A1_N(_04617_),
    .A2_N(_04604_),
    .B1(_04599_),
    .B2(_04605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_2 _13823_ (.A(\b_l[4] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04730_));
 sky130_fd_sc_hd__nand2_2 _13824_ (.A(\b_l[3] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04731_));
 sky130_fd_sc_hd__nand2_2 _13825_ (.A(_04730_),
    .B(_04731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04732_));
 sky130_fd_sc_hd__nand2_2 _13826_ (.A(\b_l[4] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04733_));
 sky130_fd_sc_hd__nand4_2 _13827_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_2 _13828_ (.A(\b_l[5] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04735_));
 sky130_fd_sc_hd__a22oi_2 _13829_ (.A1(\b_l[5] ),
    .A2(\a_h[7] ),
    .B1(_04732_),
    .B2(_04734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04736_));
 sky130_fd_sc_hd__and4_2 _13830_ (.A(_04732_),
    .B(_04734_),
    .C(\b_l[5] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04737_));
 sky130_fd_sc_hd__and3_2 _13831_ (.A(_04732_),
    .B(_04734_),
    .C(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04738_));
 sky130_fd_sc_hd__a21oi_2 _13832_ (.A1(_04732_),
    .A2(_04734_),
    .B1(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04739_));
 sky130_fd_sc_hd__nor2_2 _13833_ (.A(_04736_),
    .B(_04737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04740_));
 sky130_fd_sc_hd__nor2_2 _13834_ (.A(_04738_),
    .B(_04739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04741_));
 sky130_fd_sc_hd__o21ai_2 _13835_ (.A1(_04592_),
    .A2(_04595_),
    .B1(_04597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_2 _13836_ (.A(\b_l[2] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_2 _13837_ (.A(\b_l[1] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_2 _13838_ (.A(\b_l[0] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04745_));
 sky130_fd_sc_hd__a22oi_2 _13839_ (.A1(\b_l[1] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04746_));
 sky130_fd_sc_hd__nand2_2 _13840_ (.A(_04744_),
    .B(_04745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04747_));
 sky130_fd_sc_hd__nor2_2 _13841_ (.A(_02502_),
    .B(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04748_));
 sky130_fd_sc_hd__nand4_2 _13842_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04749_));
 sky130_fd_sc_hd__o21ai_2 _13843_ (.A1(_04746_),
    .A2(_04748_),
    .B1(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04750_));
 sky130_fd_sc_hd__o2111ai_2 _13844_ (.A1(_02502_),
    .A2(_04134_),
    .B1(\b_l[2] ),
    .C1(\a_h[10] ),
    .D1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04751_));
 sky130_fd_sc_hd__a21oi_2 _13845_ (.A1(_04747_),
    .A2(_04749_),
    .B1(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04752_));
 sky130_fd_sc_hd__o211ai_2 _13846_ (.A1(_02502_),
    .A2(_04134_),
    .B1(_04743_),
    .C1(_04747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04753_));
 sky130_fd_sc_hd__o211ai_2 _13847_ (.A1(_04592_),
    .A2(_04595_),
    .B1(_04597_),
    .C1(_04753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04754_));
 sky130_fd_sc_hd__a21oi_2 _13848_ (.A1(_04750_),
    .A2(_04751_),
    .B1(_04742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04755_));
 sky130_fd_sc_hd__nand3_2 _13849_ (.A(_04750_),
    .B(_04751_),
    .C(_04742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04756_));
 sky130_fd_sc_hd__inv_2 _13850_ (.A(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04757_));
 sky130_fd_sc_hd__o21ai_2 _13851_ (.A1(_04752_),
    .A2(_04754_),
    .B1(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_2 _13852_ (.A(_04758_),
    .B(_04740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04759_));
 sky130_fd_sc_hd__o22ai_2 _13853_ (.A1(_04736_),
    .A2(_04737_),
    .B1(_04752_),
    .B2(_04754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04760_));
 sky130_fd_sc_hd__o211ai_2 _13854_ (.A1(_04752_),
    .A2(_04754_),
    .B1(_04756_),
    .C1(_04740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04761_));
 sky130_fd_sc_hd__inv_2 _13855_ (.A(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04762_));
 sky130_fd_sc_hd__o21ai_2 _13856_ (.A1(_04736_),
    .A2(_04737_),
    .B1(_04758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04763_));
 sky130_fd_sc_hd__a21o_2 _13857_ (.A1(_04741_),
    .A2(_04758_),
    .B1(_04729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04764_));
 sky130_fd_sc_hd__and3_2 _13858_ (.A(_04763_),
    .B(_04728_),
    .C(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04765_));
 sky130_fd_sc_hd__nand3_2 _13859_ (.A(_04763_),
    .B(_04728_),
    .C(_04761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04766_));
 sky130_fd_sc_hd__o211ai_2 _13860_ (.A1(_04760_),
    .A2(_04757_),
    .B1(_04729_),
    .C1(_04759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04767_));
 sky130_fd_sc_hd__inv_2 _13861_ (.A(_04767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04768_));
 sky130_fd_sc_hd__nand2_2 _13862_ (.A(_04766_),
    .B(_04767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04769_));
 sky130_fd_sc_hd__o21ai_2 _13863_ (.A1(_04723_),
    .A2(_04726_),
    .B1(_04767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04770_));
 sky130_fd_sc_hd__a21o_2 _13864_ (.A1(_04766_),
    .A2(_04767_),
    .B1(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04771_));
 sky130_fd_sc_hd__o2111ai_2 _13865_ (.A1(_04725_),
    .A2(_04718_),
    .B1(_04724_),
    .C1(_04766_),
    .D1(_04767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04772_));
 sky130_fd_sc_hd__o21ai_2 _13866_ (.A1(_04723_),
    .A2(_04726_),
    .B1(_04769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04773_));
 sky130_fd_sc_hd__nand3_2 _13867_ (.A(_04773_),
    .B(_04652_),
    .C(_04772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04774_));
 sky130_fd_sc_hd__o211a_2 _13868_ (.A1(_04770_),
    .A2(_04765_),
    .B1(_04653_),
    .C1(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04775_));
 sky130_fd_sc_hd__o211ai_2 _13869_ (.A1(_04770_),
    .A2(_04765_),
    .B1(_04653_),
    .C1(_04771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04776_));
 sky130_fd_sc_hd__a32oi_2 _13870_ (.A1(_04629_),
    .A2(_04639_),
    .A3(_04640_),
    .B1(_04641_),
    .B2(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04777_));
 sky130_fd_sc_hd__a32o_2 _13871_ (.A1(_04629_),
    .A2(_04639_),
    .A3(_04640_),
    .B1(_04641_),
    .B2(_04627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04778_));
 sky130_fd_sc_hd__nand2_2 _13872_ (.A(\b_l[11] ),
    .B(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04779_));
 sky130_fd_sc_hd__nand2_2 _13873_ (.A(\b_l[10] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_2 _13874_ (.A(\b_l[9] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04781_));
 sky130_fd_sc_hd__a22oi_2 _13875_ (.A1(\b_l[10] ),
    .A2(\a_h[2] ),
    .B1(\a_h[3] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04782_));
 sky130_fd_sc_hd__nand2_2 _13876_ (.A(_04780_),
    .B(_04781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04783_));
 sky130_fd_sc_hd__nand4_2 _13877_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04784_));
 sky130_fd_sc_hd__nand4_2 _13878_ (.A(_04783_),
    .B(_04784_),
    .C(\b_l[11] ),
    .D(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04785_));
 sky130_fd_sc_hd__a22o_2 _13879_ (.A1(\b_l[11] ),
    .A2(\a_h[1] ),
    .B1(_04783_),
    .B2(_04784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04786_));
 sky130_fd_sc_hd__a21oi_2 _13880_ (.A1(_04661_),
    .A2(_04664_),
    .B1(_04662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04787_));
 sky130_fd_sc_hd__nand3_2 _13881_ (.A(_04785_),
    .B(_04786_),
    .C(_04787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04788_));
 sky130_fd_sc_hd__nand3_2 _13882_ (.A(_04779_),
    .B(_04783_),
    .C(_04784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04789_));
 sky130_fd_sc_hd__a21o_2 _13883_ (.A1(_04783_),
    .A2(_04784_),
    .B1(_04779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04790_));
 sky130_fd_sc_hd__nand3b_2 _13884_ (.A_N(_04787_),
    .B(_04789_),
    .C(_04790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_2 _13885_ (.A(_09177_),
    .B(_09329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04792_));
 sky130_fd_sc_hd__o211ai_2 _13886_ (.A1(_09177_),
    .A2(_09329_),
    .B1(_04788_),
    .C1(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04793_));
 sky130_fd_sc_hd__a21bo_2 _13887_ (.A1(_04788_),
    .A2(_04791_),
    .B1_N(_04792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04794_));
 sky130_fd_sc_hd__a22o_2 _13888_ (.A1(\a_h[0] ),
    .A2(\b_l[12] ),
    .B1(_04788_),
    .B2(_04791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04795_));
 sky130_fd_sc_hd__nand4_2 _13889_ (.A(_04788_),
    .B(_04791_),
    .C(\a_h[0] ),
    .D(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04796_));
 sky130_fd_sc_hd__nand3_2 _13890_ (.A(_04778_),
    .B(_04793_),
    .C(_04794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04797_));
 sky130_fd_sc_hd__nand3_2 _13891_ (.A(_04795_),
    .B(_04796_),
    .C(_04777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04798_));
 sky130_fd_sc_hd__inv_2 _13892_ (.A(_04798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04799_));
 sky130_fd_sc_hd__and3_2 _13893_ (.A(_04797_),
    .B(_04798_),
    .C(_04667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04800_));
 sky130_fd_sc_hd__nand3_2 _13894_ (.A(_04797_),
    .B(_04798_),
    .C(_04667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04801_));
 sky130_fd_sc_hd__a21oi_2 _13895_ (.A1(_04797_),
    .A2(_04798_),
    .B1(_04667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_2 _13896_ (.A1(_04797_),
    .A2(_04798_),
    .B1(_04667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04803_));
 sky130_fd_sc_hd__and3_2 _13897_ (.A(_04668_),
    .B(_04797_),
    .C(_04798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04804_));
 sky130_fd_sc_hd__a21oi_2 _13898_ (.A1(_04797_),
    .A2(_04798_),
    .B1(_04668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04805_));
 sky130_fd_sc_hd__o211ai_2 _13899_ (.A1(_04800_),
    .A2(_04802_),
    .B1(_04774_),
    .C1(_04776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04806_));
 sky130_fd_sc_hd__o2bb2ai_2 _13900_ (.A1_N(_04774_),
    .A2_N(_04776_),
    .B1(_04804_),
    .B2(_04805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04807_));
 sky130_fd_sc_hd__nand3_2 _13901_ (.A(_04774_),
    .B(_04801_),
    .C(_04803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04808_));
 sky130_fd_sc_hd__nand4_2 _13902_ (.A(_04774_),
    .B(_04776_),
    .C(_04801_),
    .D(_04803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04809_));
 sky130_fd_sc_hd__o2bb2ai_2 _13903_ (.A1_N(_04774_),
    .A2_N(_04776_),
    .B1(_04800_),
    .B2(_04802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04810_));
 sky130_fd_sc_hd__nand3_2 _13904_ (.A(_04810_),
    .B(_04702_),
    .C(_04809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04811_));
 sky130_fd_sc_hd__inv_2 _13905_ (.A(_04811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04812_));
 sky130_fd_sc_hd__o211ai_2 _13906_ (.A1(_04654_),
    .A2(_04682_),
    .B1(_04806_),
    .C1(_04807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04813_));
 sky130_fd_sc_hd__nand2_2 _13907_ (.A(_04811_),
    .B(_04813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_2 _13908_ (.A(_04813_),
    .B(_04673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_2 _13909_ (.A(_04811_),
    .B(_04813_),
    .C(_04673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04816_));
 sky130_fd_sc_hd__o2bb2ai_2 _13910_ (.A1_N(_04811_),
    .A2_N(_04813_),
    .B1(_04670_),
    .B2(_04672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04817_));
 sky130_fd_sc_hd__o21ai_2 _13911_ (.A1(_04815_),
    .A2(_04812_),
    .B1(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04818_));
 sky130_fd_sc_hd__o21ai_2 _13912_ (.A1(_04670_),
    .A2(_04672_),
    .B1(_04813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_2 _13913_ (.A(_04814_),
    .B(_04673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04820_));
 sky130_fd_sc_hd__o211ai_2 _13914_ (.A1(_04819_),
    .A2(_04812_),
    .B1(_04701_),
    .C1(_04820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04821_));
 sky130_fd_sc_hd__o211a_2 _13915_ (.A1(_04680_),
    .A2(_04700_),
    .B1(_04816_),
    .C1(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04822_));
 sky130_fd_sc_hd__o211ai_2 _13916_ (.A1(_04680_),
    .A2(_04700_),
    .B1(_04816_),
    .C1(_04817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_2 _13917_ (.A(_04821_),
    .B(_04823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04824_));
 sky130_fd_sc_hd__a32oi_2 _13918_ (.A1(_04688_),
    .A2(_04689_),
    .A3(_04690_),
    .B1(_04821_),
    .B2(_04823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04825_));
 sky130_fd_sc_hd__nor2_2 _13919_ (.A(_04693_),
    .B(_04822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04826_));
 sky130_fd_sc_hd__nor2_2 _13920_ (.A(_04693_),
    .B(_04824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04827_));
 sky130_fd_sc_hd__a21oi_2 _13921_ (.A1(_04826_),
    .A2(_04821_),
    .B1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04828_));
 sky130_fd_sc_hd__a21o_2 _13922_ (.A1(_04826_),
    .A2(_04821_),
    .B1(_04825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04829_));
 sky130_fd_sc_hd__o21ai_2 _13923_ (.A1(_04579_),
    .A2(_04691_),
    .B1(_04581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04830_));
 sky130_fd_sc_hd__a21oi_2 _13924_ (.A1(_04485_),
    .A2(_04580_),
    .B1(_04830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04831_));
 sky130_fd_sc_hd__o31ai_2 _13925_ (.A1(_04694_),
    .A2(_04829_),
    .A3(_04831_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04832_));
 sky130_fd_sc_hd__a31oi_2 _13926_ (.A1(_04696_),
    .A2(_04699_),
    .A3(_04829_),
    .B1(_04832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00318_));
 sky130_fd_sc_hd__a31o_2 _13927_ (.A1(_04777_),
    .A2(_04795_),
    .A3(_04796_),
    .B1(_04800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04833_));
 sky130_fd_sc_hd__nand2_2 _13928_ (.A(_04776_),
    .B(_04808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04834_));
 sky130_fd_sc_hd__a31oi_2 _13929_ (.A1(_04774_),
    .A2(_04801_),
    .A3(_04803_),
    .B1(_04775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04835_));
 sky130_fd_sc_hd__a22oi_2 _13930_ (.A1(\a_h[0] ),
    .A2(\b_l[13] ),
    .B1(\a_h[1] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04836_));
 sky130_fd_sc_hd__or4b_2 _13931_ (.A(_09177_),
    .B(_09329_),
    .C(_09351_),
    .D_N(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04837_));
 sky130_fd_sc_hd__a31oi_2 _13932_ (.A1(\b_l[13] ),
    .A2(\a_h[1] ),
    .A3(_04792_),
    .B1(_04836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04838_));
 sky130_fd_sc_hd__a31o_2 _13933_ (.A1(\b_l[13] ),
    .A2(\a_h[1] ),
    .A3(_04792_),
    .B1(_04836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04839_));
 sky130_fd_sc_hd__o21ai_2 _13934_ (.A1(_04779_),
    .A2(_04782_),
    .B1(_04784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_2 _13935_ (.A(\b_l[10] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_2 _13936_ (.A(\b_l[9] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04842_));
 sky130_fd_sc_hd__a22oi_2 _13937_ (.A1(\b_l[10] ),
    .A2(\a_h[3] ),
    .B1(\a_h[4] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04843_));
 sky130_fd_sc_hd__nand2_2 _13938_ (.A(_04841_),
    .B(_04842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04844_));
 sky130_fd_sc_hd__nand4_2 _13939_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[3] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04845_));
 sky130_fd_sc_hd__nand2_2 _13940_ (.A(\b_l[11] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04846_));
 sky130_fd_sc_hd__o2bb2ai_2 _13941_ (.A1_N(_04844_),
    .A2_N(_04845_),
    .B1(_09308_),
    .B2(_09395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04847_));
 sky130_fd_sc_hd__o2111ai_2 _13942_ (.A1(_01888_),
    .A2(_04555_),
    .B1(\b_l[11] ),
    .C1(\a_h[2] ),
    .D1(_04844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04848_));
 sky130_fd_sc_hd__nand3_2 _13943_ (.A(_04847_),
    .B(_04848_),
    .C(_04840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04849_));
 sky130_fd_sc_hd__a21oi_2 _13944_ (.A1(_04844_),
    .A2(_04845_),
    .B1(_04846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04850_));
 sky130_fd_sc_hd__o21a_2 _13945_ (.A1(_01888_),
    .A2(_04555_),
    .B1(_04846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04851_));
 sky130_fd_sc_hd__nand2_2 _13946_ (.A(_04845_),
    .B(_04846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04852_));
 sky130_fd_sc_hd__o221ai_2 _13947_ (.A1(_04779_),
    .A2(_04782_),
    .B1(_04843_),
    .B2(_04852_),
    .C1(_04784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04853_));
 sky130_fd_sc_hd__a21o_2 _13948_ (.A1(_04847_),
    .A2(_04848_),
    .B1(_04840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04854_));
 sky130_fd_sc_hd__o21ai_2 _13949_ (.A1(_04850_),
    .A2(_04853_),
    .B1(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_2 _13950_ (.A(_04839_),
    .B(_04855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04856_));
 sky130_fd_sc_hd__o211ai_2 _13951_ (.A1(_04850_),
    .A2(_04853_),
    .B1(_04838_),
    .C1(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04857_));
 sky130_fd_sc_hd__o211ai_2 _13952_ (.A1(_04850_),
    .A2(_04853_),
    .B1(_04839_),
    .C1(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_2 _13953_ (.A(_04855_),
    .B(_04838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04859_));
 sky130_fd_sc_hd__o22ai_2 _13954_ (.A1(_04608_),
    .A2(_04720_),
    .B1(_04722_),
    .B2(_04718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04860_));
 sky130_fd_sc_hd__nand2_2 _13955_ (.A(_04719_),
    .B(_04725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04861_));
 sky130_fd_sc_hd__and3_2 _13956_ (.A(_04858_),
    .B(_04859_),
    .C(_04861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04862_));
 sky130_fd_sc_hd__nand3_2 _13957_ (.A(_04858_),
    .B(_04859_),
    .C(_04861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04863_));
 sky130_fd_sc_hd__nand3_2 _13958_ (.A(_04856_),
    .B(_04857_),
    .C(_04860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04864_));
 sky130_fd_sc_hd__nand2_2 _13959_ (.A(_04863_),
    .B(_04864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04865_));
 sky130_fd_sc_hd__a21boi_2 _13960_ (.A1(_04791_),
    .A2(_04792_),
    .B1_N(_04788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04866_));
 sky130_fd_sc_hd__a31o_2 _13961_ (.A1(_04856_),
    .A2(_04857_),
    .A3(_04860_),
    .B1(_04866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_2 _13962_ (.A(_04865_),
    .B(_04866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04868_));
 sky130_fd_sc_hd__o21ai_2 _13963_ (.A1(_04862_),
    .A2(_04867_),
    .B1(_04868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04869_));
 sky130_fd_sc_hd__a31oi_2 _13964_ (.A1(_04728_),
    .A2(_04761_),
    .A3(_04763_),
    .B1(_04727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04870_));
 sky130_fd_sc_hd__o2bb2ai_2 _13965_ (.A1_N(_04727_),
    .A2_N(_04767_),
    .B1(_04762_),
    .B2(_04764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04871_));
 sky130_fd_sc_hd__o21a_2 _13966_ (.A1(_04736_),
    .A2(_04737_),
    .B1(_04756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04872_));
 sky130_fd_sc_hd__a2bb2oi_2 _13967_ (.A1_N(_04752_),
    .A2_N(_04754_),
    .B1(_04756_),
    .B2(_04741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2_2 _13968_ (.A(\b_l[5] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_2 _13969_ (.A(\b_l[3] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04875_));
 sky130_fd_sc_hd__and4_2 _13970_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04876_));
 sky130_fd_sc_hd__nand4_2 _13971_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04877_));
 sky130_fd_sc_hd__a22oi_2 _13972_ (.A1(\b_l[4] ),
    .A2(\a_h[9] ),
    .B1(\a_h[10] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04878_));
 sky130_fd_sc_hd__nand2_2 _13973_ (.A(_04733_),
    .B(_04875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04879_));
 sky130_fd_sc_hd__o211a_2 _13974_ (.A1(_04876_),
    .A2(_04878_),
    .B1(\b_l[5] ),
    .C1(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04880_));
 sky130_fd_sc_hd__o311a_2 _13975_ (.A1(_09471_),
    .A2(_09482_),
    .A3(_04182_),
    .B1(_04874_),
    .C1(_04879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04881_));
 sky130_fd_sc_hd__a21oi_2 _13976_ (.A1(_04733_),
    .A2(_04875_),
    .B1(_04874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04882_));
 sky130_fd_sc_hd__a21o_2 _13977_ (.A1(_04733_),
    .A2(_04875_),
    .B1(_04874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04883_));
 sky130_fd_sc_hd__and4_2 _13978_ (.A(_04879_),
    .B(\a_h[8] ),
    .C(\b_l[5] ),
    .D(_04877_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04884_));
 sky130_fd_sc_hd__o22a_2 _13979_ (.A1(_09220_),
    .A2(_09460_),
    .B1(_04876_),
    .B2(_04878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04885_));
 sky130_fd_sc_hd__a22o_2 _13980_ (.A1(\b_l[5] ),
    .A2(\a_h[8] ),
    .B1(_04877_),
    .B2(_04879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04886_));
 sky130_fd_sc_hd__o21ai_2 _13981_ (.A1(_04876_),
    .A2(_04883_),
    .B1(_04886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04887_));
 sky130_fd_sc_hd__o21a_2 _13982_ (.A1(_04876_),
    .A2(_04883_),
    .B1(_04886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04888_));
 sky130_fd_sc_hd__a21oi_2 _13983_ (.A1(_04744_),
    .A2(_04745_),
    .B1(_04743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04889_));
 sky130_fd_sc_hd__o22a_2 _13984_ (.A1(_09155_),
    .A2(_09482_),
    .B1(_02502_),
    .B2(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04890_));
 sky130_fd_sc_hd__and2_2 _13985_ (.A(\b_l[2] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04891_));
 sky130_fd_sc_hd__nand2_2 _13986_ (.A(\b_l[2] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_2 _13987_ (.A(\b_l[0] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_2 _13988_ (.A(\b_l[1] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04894_));
 sky130_fd_sc_hd__a22oi_2 _13989_ (.A1(\b_l[1] ),
    .A2(\a_h[12] ),
    .B1(\a_h[13] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04895_));
 sky130_fd_sc_hd__nand2_2 _13990_ (.A(_04893_),
    .B(_04894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04896_));
 sky130_fd_sc_hd__nand3_2 _13991_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04897_));
 sky130_fd_sc_hd__nand4_2 _13992_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04898_));
 sky130_fd_sc_hd__o211a_2 _13993_ (.A1(_09515_),
    .A2(_04897_),
    .B1(_04891_),
    .C1(_04896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04899_));
 sky130_fd_sc_hd__o2111ai_2 _13994_ (.A1(_09515_),
    .A2(_04897_),
    .B1(\a_h[11] ),
    .C1(_04896_),
    .D1(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04900_));
 sky130_fd_sc_hd__a21oi_2 _13995_ (.A1(_04896_),
    .A2(_04898_),
    .B1(_04891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04901_));
 sky130_fd_sc_hd__o2bb2ai_2 _13996_ (.A1_N(_04896_),
    .A2_N(_04898_),
    .B1(_09155_),
    .B2(_09493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04902_));
 sky130_fd_sc_hd__o211a_2 _13997_ (.A1(_04748_),
    .A2(_04889_),
    .B1(_04900_),
    .C1(_04902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04903_));
 sky130_fd_sc_hd__o211ai_2 _13998_ (.A1(_04748_),
    .A2(_04889_),
    .B1(_04900_),
    .C1(_04902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04904_));
 sky130_fd_sc_hd__a2bb2oi_2 _13999_ (.A1_N(_04746_),
    .A2_N(_04890_),
    .B1(_04900_),
    .B2(_04902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04905_));
 sky130_fd_sc_hd__o22ai_2 _14000_ (.A1(_04746_),
    .A2(_04890_),
    .B1(_04899_),
    .B2(_04901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2_2 _14001_ (.A(_04904_),
    .B(_04906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04907_));
 sky130_fd_sc_hd__o211ai_2 _14002_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04904_),
    .C1(_04906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04908_));
 sky130_fd_sc_hd__inv_2 _14003_ (.A(_04908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04909_));
 sky130_fd_sc_hd__o22ai_2 _14004_ (.A1(_04880_),
    .A2(_04881_),
    .B1(_04903_),
    .B2(_04905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04910_));
 sky130_fd_sc_hd__nand3_2 _14005_ (.A(_04888_),
    .B(_04904_),
    .C(_04906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04911_));
 sky130_fd_sc_hd__o22ai_2 _14006_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04903_),
    .B2(_04905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04912_));
 sky130_fd_sc_hd__nand3_2 _14007_ (.A(_04912_),
    .B(_04873_),
    .C(_04911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04913_));
 sky130_fd_sc_hd__a21oi_2 _14008_ (.A1(_04888_),
    .A2(_04907_),
    .B1(_04873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04914_));
 sky130_fd_sc_hd__o21ai_2 _14009_ (.A1(_04755_),
    .A2(_04872_),
    .B1(_04910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04915_));
 sky130_fd_sc_hd__o211ai_2 _14010_ (.A1(_04755_),
    .A2(_04872_),
    .B1(_04908_),
    .C1(_04910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_2 _14011_ (.A(_04913_),
    .B(_04916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04917_));
 sky130_fd_sc_hd__a31o_2 _14012_ (.A1(\b_l[8] ),
    .A2(_04711_),
    .A3(\a_h[4] ),
    .B1(_04709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04918_));
 sky130_fd_sc_hd__nand2_2 _14013_ (.A(_04734_),
    .B(_04735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_2 _14014_ (.A(_04732_),
    .B(_04919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04920_));
 sky130_fd_sc_hd__a21boi_2 _14015_ (.A1(_04734_),
    .A2(_04735_),
    .B1_N(_04732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_2 _14016_ (.A(\b_l[8] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_2 _14017_ (.A(\b_l[6] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04923_));
 sky130_fd_sc_hd__a22o_2 _14018_ (.A1(\b_l[7] ),
    .A2(\a_h[6] ),
    .B1(\a_h[7] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04924_));
 sky130_fd_sc_hd__nand2_2 _14019_ (.A(\b_l[7] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04925_));
 sky130_fd_sc_hd__nand4_2 _14020_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[6] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04926_));
 sky130_fd_sc_hd__o2bb2ai_2 _14021_ (.A1_N(_04707_),
    .A2_N(_04923_),
    .B1(_04925_),
    .B2(_04708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04927_));
 sky130_fd_sc_hd__o2111ai_2 _14022_ (.A1(_04708_),
    .A2(_04925_),
    .B1(\b_l[8] ),
    .C1(\a_h[5] ),
    .D1(_04924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04928_));
 sky130_fd_sc_hd__o21ai_2 _14023_ (.A1(_09264_),
    .A2(_09428_),
    .B1(_04927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04929_));
 sky130_fd_sc_hd__o221ai_2 _14024_ (.A1(_09264_),
    .A2(_09428_),
    .B1(_04708_),
    .B2(_04925_),
    .C1(_04924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04930_));
 sky130_fd_sc_hd__nand3_2 _14025_ (.A(_04927_),
    .B(\a_h[5] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04931_));
 sky130_fd_sc_hd__nand3_2 _14026_ (.A(_04921_),
    .B(_04928_),
    .C(_04929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04932_));
 sky130_fd_sc_hd__nand3_2 _14027_ (.A(_04931_),
    .B(_04920_),
    .C(_04930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04933_));
 sky130_fd_sc_hd__and2_2 _14028_ (.A(_04933_),
    .B(_04918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04934_));
 sky130_fd_sc_hd__nand2_2 _14029_ (.A(_04933_),
    .B(_04918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04935_));
 sky130_fd_sc_hd__and3_2 _14030_ (.A(_04932_),
    .B(_04933_),
    .C(_04918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04936_));
 sky130_fd_sc_hd__a21oi_2 _14031_ (.A1(_04932_),
    .A2(_04933_),
    .B1(_04918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04937_));
 sky130_fd_sc_hd__a21oi_2 _14032_ (.A1(_04934_),
    .A2(_04932_),
    .B1(_04937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04938_));
 sky130_fd_sc_hd__a21o_2 _14033_ (.A1(_04934_),
    .A2(_04932_),
    .B1(_04937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04939_));
 sky130_fd_sc_hd__o221a_2 _14034_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04909_),
    .B2(_04915_),
    .C1(_04913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04940_));
 sky130_fd_sc_hd__o221ai_2 _14035_ (.A1(_04936_),
    .A2(_04937_),
    .B1(_04909_),
    .B2(_04915_),
    .C1(_04913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04941_));
 sky130_fd_sc_hd__a21o_2 _14036_ (.A1(_04913_),
    .A2(_04916_),
    .B1(_04939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04942_));
 sky130_fd_sc_hd__nand3_2 _14037_ (.A(_04913_),
    .B(_04916_),
    .C(_04938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04943_));
 sky130_fd_sc_hd__o2bb2ai_2 _14038_ (.A1_N(_04913_),
    .A2_N(_04916_),
    .B1(_04936_),
    .B2(_04937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04944_));
 sky130_fd_sc_hd__nand3_2 _14039_ (.A(_04944_),
    .B(_04871_),
    .C(_04943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04945_));
 sky130_fd_sc_hd__o2bb2ai_2 _14040_ (.A1_N(_04917_),
    .A2_N(_04938_),
    .B1(_04768_),
    .B2(_04870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04946_));
 sky130_fd_sc_hd__o211ai_2 _14041_ (.A1(_04768_),
    .A2(_04870_),
    .B1(_04941_),
    .C1(_04942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04947_));
 sky130_fd_sc_hd__o211ai_2 _14042_ (.A1(_04940_),
    .A2(_04946_),
    .B1(_04945_),
    .C1(_04869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04948_));
 sky130_fd_sc_hd__a21o_2 _14043_ (.A1(_04945_),
    .A2(_04947_),
    .B1(_04869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04949_));
 sky130_fd_sc_hd__a21bo_2 _14044_ (.A1(_04945_),
    .A2(_04947_),
    .B1_N(_04869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04950_));
 sky130_fd_sc_hd__o2111ai_2 _14045_ (.A1(_04862_),
    .A2(_04867_),
    .B1(_04868_),
    .C1(_04945_),
    .D1(_04947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04951_));
 sky130_fd_sc_hd__nand3_2 _14046_ (.A(_04835_),
    .B(_04948_),
    .C(_04949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04952_));
 sky130_fd_sc_hd__nand3_2 _14047_ (.A(_04950_),
    .B(_04951_),
    .C(_04834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04953_));
 sky130_fd_sc_hd__a21oi_2 _14048_ (.A1(_04952_),
    .A2(_04953_),
    .B1(_04833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04954_));
 sky130_fd_sc_hd__a21o_2 _14049_ (.A1(_04952_),
    .A2(_04953_),
    .B1(_04833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04955_));
 sky130_fd_sc_hd__o211a_2 _14050_ (.A1(_04799_),
    .A2(_04800_),
    .B1(_04952_),
    .C1(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04956_));
 sky130_fd_sc_hd__o211ai_2 _14051_ (.A1(_04799_),
    .A2(_04800_),
    .B1(_04952_),
    .C1(_04953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04957_));
 sky130_fd_sc_hd__nand2_2 _14052_ (.A(_04811_),
    .B(_04815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04958_));
 sky130_fd_sc_hd__o21bai_2 _14053_ (.A1(_04954_),
    .A2(_04956_),
    .B1_N(_04958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04959_));
 sky130_fd_sc_hd__and3_2 _14054_ (.A(_04955_),
    .B(_04957_),
    .C(_04958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04960_));
 sky130_fd_sc_hd__nand3_2 _14055_ (.A(_04955_),
    .B(_04957_),
    .C(_04958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04961_));
 sky130_fd_sc_hd__o2bb2ai_2 _14056_ (.A1_N(_04959_),
    .A2_N(_04961_),
    .B1(_04701_),
    .B2(_04818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04962_));
 sky130_fd_sc_hd__nand3_2 _14057_ (.A(_04959_),
    .B(_04961_),
    .C(_04822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_2 _14058_ (.A(_04962_),
    .B(_04963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04964_));
 sky130_fd_sc_hd__o32a_2 _14059_ (.A1(_04694_),
    .A2(_04829_),
    .A3(_04831_),
    .B1(_04824_),
    .B2(_04693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04965_));
 sky130_fd_sc_hd__o21ai_2 _14060_ (.A1(_04964_),
    .A2(_04965_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_2 _14061_ (.A1(_04964_),
    .A2(_04965_),
    .B1(_04966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00319_));
 sky130_fd_sc_hd__o2bb2ai_2 _14062_ (.A1_N(_04869_),
    .A2_N(_04945_),
    .B1(_04940_),
    .B2(_04946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04967_));
 sky130_fd_sc_hd__o2bb2ai_2 _14063_ (.A1_N(_04913_),
    .A2_N(_04939_),
    .B1(_04915_),
    .B2(_04909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04968_));
 sky130_fd_sc_hd__a22oi_2 _14064_ (.A1(_04914_),
    .A2(_04908_),
    .B1(_04913_),
    .B2(_04939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04969_));
 sky130_fd_sc_hd__o21ai_2 _14065_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04970_));
 sky130_fd_sc_hd__o21ai_2 _14066_ (.A1(_04887_),
    .A2(_04905_),
    .B1(_04904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_2 _14067_ (.A(_04906_),
    .B(_04970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_2 _14068_ (.A(\b_l[5] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04973_));
 sky130_fd_sc_hd__a22oi_2 _14069_ (.A1(\b_l[4] ),
    .A2(\a_h[10] ),
    .B1(\a_h[11] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04974_));
 sky130_fd_sc_hd__and4_2 _14070_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04975_));
 sky130_fd_sc_hd__nand4_2 _14071_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_2 _14072_ (.A1(_02362_),
    .A2(_04182_),
    .B1(_04973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04977_));
 sky130_fd_sc_hd__o21bai_2 _14073_ (.A1(_04974_),
    .A2(_04975_),
    .B1_N(_04973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04978_));
 sky130_fd_sc_hd__o21ai_2 _14074_ (.A1(_04974_),
    .A2(_04977_),
    .B1(_04978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04979_));
 sky130_fd_sc_hd__a21o_2 _14075_ (.A1(_04892_),
    .A2(_04898_),
    .B1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04980_));
 sky130_fd_sc_hd__a21oi_2 _14076_ (.A1(_04892_),
    .A2(_04898_),
    .B1(_04895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_2 _14077_ (.A(\b_l[2] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04982_));
 sky130_fd_sc_hd__nand2_2 _14078_ (.A(\b_l[0] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_2 _14079_ (.A(\b_l[1] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04984_));
 sky130_fd_sc_hd__a22oi_2 _14080_ (.A1(\b_l[1] ),
    .A2(\a_h[13] ),
    .B1(\a_h[14] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_2 _14081_ (.A(_04983_),
    .B(_04984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04986_));
 sky130_fd_sc_hd__and2_2 _14082_ (.A(\b_l[1] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04987_));
 sky130_fd_sc_hd__nand2_2 _14083_ (.A(\b_l[1] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04988_));
 sky130_fd_sc_hd__nand4_2 _14084_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[13] ),
    .D(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04989_));
 sky130_fd_sc_hd__a22oi_2 _14085_ (.A1(\b_l[2] ),
    .A2(\a_h[12] ),
    .B1(_04986_),
    .B2(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04990_));
 sky130_fd_sc_hd__a22o_2 _14086_ (.A1(\b_l[2] ),
    .A2(\a_h[12] ),
    .B1(_04986_),
    .B2(_04989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04991_));
 sky130_fd_sc_hd__nand4_2 _14087_ (.A(_04986_),
    .B(_04989_),
    .C(\b_l[2] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_2 _14088_ (.A(_04981_),
    .B(_04992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04993_));
 sky130_fd_sc_hd__nand3_2 _14089_ (.A(_04981_),
    .B(_04991_),
    .C(_04992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04994_));
 sky130_fd_sc_hd__o221ai_2 _14090_ (.A1(_09155_),
    .A2(_09504_),
    .B1(_04893_),
    .B2(_04988_),
    .C1(_04986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04995_));
 sky130_fd_sc_hd__a21o_2 _14091_ (.A1(_04986_),
    .A2(_04989_),
    .B1(_04982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_04996_));
 sky130_fd_sc_hd__nand3_2 _14092_ (.A(_04996_),
    .B(_04980_),
    .C(_04995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04997_));
 sky130_fd_sc_hd__o21ai_2 _14093_ (.A1(_04990_),
    .A2(_04993_),
    .B1(_04997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04998_));
 sky130_fd_sc_hd__o211ai_2 _14094_ (.A1(_04990_),
    .A2(_04993_),
    .B1(_04997_),
    .C1(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_04999_));
 sky130_fd_sc_hd__o211a_2 _14095_ (.A1(_04974_),
    .A2(_04977_),
    .B1(_04978_),
    .C1(_04998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05000_));
 sky130_fd_sc_hd__a21o_2 _14096_ (.A1(_04994_),
    .A2(_04997_),
    .B1(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05001_));
 sky130_fd_sc_hd__o2111ai_2 _14097_ (.A1(_04974_),
    .A2(_04977_),
    .B1(_04978_),
    .C1(_04994_),
    .D1(_04997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05002_));
 sky130_fd_sc_hd__nand2_2 _14098_ (.A(_04998_),
    .B(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05003_));
 sky130_fd_sc_hd__nand3_2 _14099_ (.A(_04972_),
    .B(_05002_),
    .C(_05003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_2 _14100_ (.A(_04971_),
    .B(_04999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05005_));
 sky130_fd_sc_hd__nand3_2 _14101_ (.A(_05001_),
    .B(_04971_),
    .C(_04999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05006_));
 sky130_fd_sc_hd__a22o_2 _14102_ (.A1(_04707_),
    .A2(_04923_),
    .B1(_04926_),
    .B2(_04922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05007_));
 sky130_fd_sc_hd__a22oi_2 _14103_ (.A1(_04707_),
    .A2(_04923_),
    .B1(_04926_),
    .B2(_04922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05008_));
 sky130_fd_sc_hd__a21o_2 _14104_ (.A1(_04874_),
    .A2(_04877_),
    .B1(_04878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05009_));
 sky130_fd_sc_hd__and2_2 _14105_ (.A(\b_l[8] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05010_));
 sky130_fd_sc_hd__nand2_2 _14106_ (.A(\b_l[8] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05011_));
 sky130_fd_sc_hd__nand2_2 _14107_ (.A(\b_l[6] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_2 _14108_ (.A(_04925_),
    .B(_05012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05013_));
 sky130_fd_sc_hd__nand4_2 _14109_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05014_));
 sky130_fd_sc_hd__nand4_2 _14110_ (.A(_05013_),
    .B(_05014_),
    .C(\b_l[8] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05015_));
 sky130_fd_sc_hd__a21o_2 _14111_ (.A1(_05013_),
    .A2(_05014_),
    .B1(_05010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05016_));
 sky130_fd_sc_hd__a21o_2 _14112_ (.A1(_05013_),
    .A2(_05014_),
    .B1(_05011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05017_));
 sky130_fd_sc_hd__o211ai_2 _14113_ (.A1(_09264_),
    .A2(_09439_),
    .B1(_05013_),
    .C1(_05014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05018_));
 sky130_fd_sc_hd__o211ai_2 _14114_ (.A1(_04876_),
    .A2(_04882_),
    .B1(_05015_),
    .C1(_05016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05019_));
 sky130_fd_sc_hd__and3_2 _14115_ (.A(_05017_),
    .B(_05018_),
    .C(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05020_));
 sky130_fd_sc_hd__nand3_2 _14116_ (.A(_05017_),
    .B(_05018_),
    .C(_05009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_2 _14117_ (.A(_05019_),
    .B(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05022_));
 sky130_fd_sc_hd__a32oi_2 _14118_ (.A1(_05009_),
    .A2(_05017_),
    .A3(_05018_),
    .B1(_05019_),
    .B2(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_2 _14119_ (.A(_05021_),
    .B(_05022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05024_));
 sky130_fd_sc_hd__and3_2 _14120_ (.A(_05008_),
    .B(_05019_),
    .C(_05021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05025_));
 sky130_fd_sc_hd__a21oi_2 _14121_ (.A1(_05019_),
    .A2(_05021_),
    .B1(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05026_));
 sky130_fd_sc_hd__a21o_2 _14122_ (.A1(_05019_),
    .A2(_05021_),
    .B1(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05027_));
 sky130_fd_sc_hd__and3_2 _14123_ (.A(_05019_),
    .B(_05021_),
    .C(_05007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05028_));
 sky130_fd_sc_hd__a21oi_2 _14124_ (.A1(_05019_),
    .A2(_05021_),
    .B1(_05008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05029_));
 sky130_fd_sc_hd__o21ai_2 _14125_ (.A1(_05020_),
    .A2(_05022_),
    .B1(_05027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05030_));
 sky130_fd_sc_hd__nand3b_2 _14126_ (.A_N(_05030_),
    .B(_05006_),
    .C(_05004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05031_));
 sky130_fd_sc_hd__nand2_2 _14127_ (.A(_05004_),
    .B(_05030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05032_));
 sky130_fd_sc_hd__o21ai_2 _14128_ (.A1(_05000_),
    .A2(_05005_),
    .B1(_05032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05033_));
 sky130_fd_sc_hd__a21boi_2 _14129_ (.A1(_05004_),
    .A2(_05030_),
    .B1_N(_05006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05034_));
 sky130_fd_sc_hd__o211ai_2 _14130_ (.A1(_05000_),
    .A2(_05005_),
    .B1(_05030_),
    .C1(_05004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05035_));
 sky130_fd_sc_hd__o2bb2ai_2 _14131_ (.A1_N(_05004_),
    .A2_N(_05006_),
    .B1(_05026_),
    .B2(_05028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05036_));
 sky130_fd_sc_hd__nand3_2 _14132_ (.A(_04968_),
    .B(_05031_),
    .C(_05036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05037_));
 sky130_fd_sc_hd__o2bb2ai_2 _14133_ (.A1_N(_05004_),
    .A2_N(_05006_),
    .B1(_05025_),
    .B2(_05029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05038_));
 sky130_fd_sc_hd__nand3_2 _14134_ (.A(_04969_),
    .B(_05035_),
    .C(_05038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05039_));
 sky130_fd_sc_hd__a32oi_2 _14135_ (.A1(_04921_),
    .A2(_04928_),
    .A3(_04929_),
    .B1(_04933_),
    .B2(_04918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_2 _14136_ (.A(_04932_),
    .B(_04935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05041_));
 sky130_fd_sc_hd__a22oi_2 _14137_ (.A1(\b_l[13] ),
    .A2(\a_h[1] ),
    .B1(\a_h[2] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05042_));
 sky130_fd_sc_hd__and2_2 _14138_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05043_));
 sky130_fd_sc_hd__nand2_2 _14139_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05044_));
 sky130_fd_sc_hd__and4_2 _14140_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05045_));
 sky130_fd_sc_hd__nand4_2 _14141_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[1] ),
    .D(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2_2 _14142_ (.A(\a_h[0] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05047_));
 sky130_fd_sc_hd__nand3b_2 _14143_ (.A_N(_05042_),
    .B(_05046_),
    .C(_05047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05048_));
 sky130_fd_sc_hd__o21bai_2 _14144_ (.A1(_05042_),
    .A2(_05045_),
    .B1_N(_05047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_2 _14145_ (.A(_05048_),
    .B(_05049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05050_));
 sky130_fd_sc_hd__o21ai_2 _14146_ (.A1(_04846_),
    .A2(_04843_),
    .B1(_04845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_2 _14147_ (.A(\b_l[11] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05052_));
 sky130_fd_sc_hd__nand2_2 _14148_ (.A(\b_l[9] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05053_));
 sky130_fd_sc_hd__nand2_2 _14149_ (.A(\b_l[10] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_2 _14150_ (.A(_05053_),
    .B(_05054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_2 _14151_ (.A(\b_l[10] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05056_));
 sky130_fd_sc_hd__and4_2 _14152_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05057_));
 sky130_fd_sc_hd__nand4_2 _14153_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05058_));
 sky130_fd_sc_hd__o2bb2ai_2 _14154_ (.A1_N(_05055_),
    .A2_N(_05058_),
    .B1(_09308_),
    .B2(_09406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05059_));
 sky130_fd_sc_hd__o2111ai_2 _14155_ (.A1(_04842_),
    .A2(_05056_),
    .B1(\b_l[11] ),
    .C1(\a_h[3] ),
    .D1(_05055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05060_));
 sky130_fd_sc_hd__o221ai_2 _14156_ (.A1(_09308_),
    .A2(_09406_),
    .B1(_04842_),
    .B2(_05056_),
    .C1(_05055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05061_));
 sky130_fd_sc_hd__a21o_2 _14157_ (.A1(_05055_),
    .A2(_05058_),
    .B1(_05052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05062_));
 sky130_fd_sc_hd__o211ai_2 _14158_ (.A1(_04843_),
    .A2(_04851_),
    .B1(_05061_),
    .C1(_05062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05063_));
 sky130_fd_sc_hd__inv_2 _14159_ (.A(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05064_));
 sky130_fd_sc_hd__and3_2 _14160_ (.A(_05059_),
    .B(_05060_),
    .C(_05051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05065_));
 sky130_fd_sc_hd__nand3_2 _14161_ (.A(_05059_),
    .B(_05060_),
    .C(_05051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05066_));
 sky130_fd_sc_hd__nand2_2 _14162_ (.A(_05063_),
    .B(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_2 _14163_ (.A(_05067_),
    .B(_05050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05068_));
 sky130_fd_sc_hd__nand4_2 _14164_ (.A(_05048_),
    .B(_05049_),
    .C(_05063_),
    .D(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_2 _14165_ (.A(_05050_),
    .B(_05066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05070_));
 sky130_fd_sc_hd__a21o_2 _14166_ (.A1(_05063_),
    .A2(_05066_),
    .B1(_05050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05071_));
 sky130_fd_sc_hd__o211a_2 _14167_ (.A1(_05070_),
    .A2(_05064_),
    .B1(_05041_),
    .C1(_05071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05072_));
 sky130_fd_sc_hd__o211ai_2 _14168_ (.A1(_05070_),
    .A2(_05064_),
    .B1(_05041_),
    .C1(_05071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05073_));
 sky130_fd_sc_hd__nand3_2 _14169_ (.A(_05068_),
    .B(_05069_),
    .C(_05040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05074_));
 sky130_fd_sc_hd__nand2_2 _14170_ (.A(_05073_),
    .B(_05074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05075_));
 sky130_fd_sc_hd__a21boi_2 _14171_ (.A1(_04854_),
    .A2(_04838_),
    .B1_N(_04849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05076_));
 sky130_fd_sc_hd__a21oi_2 _14172_ (.A1(_05073_),
    .A2(_05074_),
    .B1(_05076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05077_));
 sky130_fd_sc_hd__and3_2 _14173_ (.A(_05073_),
    .B(_05074_),
    .C(_05076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05078_));
 sky130_fd_sc_hd__nand2_2 _14174_ (.A(_05075_),
    .B(_05076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05079_));
 sky130_fd_sc_hd__a31o_2 _14175_ (.A1(_05068_),
    .A2(_05069_),
    .A3(_05040_),
    .B1(_05076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05080_));
 sky130_fd_sc_hd__o21ai_2 _14176_ (.A1(_05072_),
    .A2(_05080_),
    .B1(_05079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05081_));
 sky130_fd_sc_hd__nand3_2 _14177_ (.A(_05037_),
    .B(_05039_),
    .C(_05081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05082_));
 sky130_fd_sc_hd__o2bb2ai_2 _14178_ (.A1_N(_05037_),
    .A2_N(_05039_),
    .B1(_05077_),
    .B2(_05078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05083_));
 sky130_fd_sc_hd__nand3_2 _14179_ (.A(_05083_),
    .B(_04967_),
    .C(_05082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05084_));
 sky130_fd_sc_hd__a21oi_2 _14180_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05085_));
 sky130_fd_sc_hd__a21o_2 _14181_ (.A1(_05082_),
    .A2(_05083_),
    .B1(_04967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05086_));
 sky130_fd_sc_hd__a21o_2 _14182_ (.A1(_04864_),
    .A2(_04866_),
    .B1(_04862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05087_));
 sky130_fd_sc_hd__and4b_2 _14183_ (.A_N(_05087_),
    .B(_04792_),
    .C(\a_h[1] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05088_));
 sky130_fd_sc_hd__inv_2 _14184_ (.A(_05088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05089_));
 sky130_fd_sc_hd__xor2_2 _14185_ (.A(_04837_),
    .B(_05087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05090_));
 sky130_fd_sc_hd__inv_2 _14186_ (.A(_05090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05091_));
 sky130_fd_sc_hd__nand2_2 _14187_ (.A(_05084_),
    .B(_05090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05092_));
 sky130_fd_sc_hd__a21o_2 _14188_ (.A1(_05084_),
    .A2(_05086_),
    .B1(_05091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05093_));
 sky130_fd_sc_hd__nand3_2 _14189_ (.A(_05084_),
    .B(_05086_),
    .C(_05091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05094_));
 sky130_fd_sc_hd__nand4_2 _14190_ (.A(_04953_),
    .B(_04957_),
    .C(_05093_),
    .D(_05094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05095_));
 sky130_fd_sc_hd__a22oi_2 _14191_ (.A1(_04953_),
    .A2(_04957_),
    .B1(_05093_),
    .B2(_05094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05096_));
 sky130_fd_sc_hd__a22o_2 _14192_ (.A1(_04953_),
    .A2(_04957_),
    .B1(_05093_),
    .B2(_05094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05097_));
 sky130_fd_sc_hd__a21oi_2 _14193_ (.A1(_05095_),
    .A2(_05097_),
    .B1(_04960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05098_));
 sky130_fd_sc_hd__a32o_2 _14194_ (.A1(_04955_),
    .A2(_04958_),
    .A3(_04957_),
    .B1(_05097_),
    .B2(_05095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05099_));
 sky130_fd_sc_hd__nand3_2 _14195_ (.A(_05097_),
    .B(_04960_),
    .C(_05095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05100_));
 sky130_fd_sc_hd__a32oi_2 _14196_ (.A1(_04822_),
    .A2(_04959_),
    .A3(_04961_),
    .B1(_04962_),
    .B2(_04827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05101_));
 sky130_fd_sc_hd__nand4_2 _14197_ (.A(_04828_),
    .B(_04962_),
    .C(_04963_),
    .D(_04695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05102_));
 sky130_fd_sc_hd__o41a_2 _14198_ (.A1(_04694_),
    .A2(_04829_),
    .A3(_04964_),
    .A4(_04831_),
    .B1(_05101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05103_));
 sky130_fd_sc_hd__a21bo_2 _14199_ (.A1(_05099_),
    .A2(_05100_),
    .B1_N(_05103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05104_));
 sky130_fd_sc_hd__or3b_2 _14200_ (.A(_05098_),
    .B(_05103_),
    .C_N(_05100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05105_));
 sky130_fd_sc_hd__and3_2 _14201_ (.A(_09690_),
    .B(_05104_),
    .C(_05105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00320_));
 sky130_fd_sc_hd__nand2_2 _14202_ (.A(_05086_),
    .B(_05092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05106_));
 sky130_fd_sc_hd__a21oi_2 _14203_ (.A1(_05084_),
    .A2(_05090_),
    .B1(_05085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05107_));
 sky130_fd_sc_hd__o32a_2 _14204_ (.A1(_09329_),
    .A2(_09351_),
    .A3(_01860_),
    .B1(_05042_),
    .B2(_05047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05108_));
 sky130_fd_sc_hd__a21o_2 _14205_ (.A1(_05073_),
    .A2(_05080_),
    .B1(_05108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05109_));
 sky130_fd_sc_hd__inv_2 _14206_ (.A(_05109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05110_));
 sky130_fd_sc_hd__and3_2 _14207_ (.A(_05073_),
    .B(_05080_),
    .C(_05108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05111_));
 sky130_fd_sc_hd__nand3_2 _14208_ (.A(_05073_),
    .B(_05080_),
    .C(_05108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05112_));
 sky130_fd_sc_hd__o21a_2 _14209_ (.A1(_09177_),
    .A2(_09384_),
    .B1(_05109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05113_));
 sky130_fd_sc_hd__a22o_2 _14210_ (.A1(\a_h[0] ),
    .A2(\b_l[15] ),
    .B1(_05109_),
    .B2(_05112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05114_));
 sky130_fd_sc_hd__nand4_2 _14211_ (.A(_05109_),
    .B(_05112_),
    .C(\a_h[0] ),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_2 _14212_ (.A(_05114_),
    .B(_05115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05116_));
 sky130_fd_sc_hd__nand2_2 _14213_ (.A(_05039_),
    .B(_05081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05117_));
 sky130_fd_sc_hd__a32oi_2 _14214_ (.A1(_04968_),
    .A2(_05031_),
    .A3(_05036_),
    .B1(_05039_),
    .B2(_05081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_2 _14215_ (.A(_05037_),
    .B(_05117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05119_));
 sky130_fd_sc_hd__a32o_2 _14216_ (.A1(\a_h[7] ),
    .A2(\a_h[8] ),
    .A3(_04259_),
    .B1(_05010_),
    .B2(_05013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05120_));
 sky130_fd_sc_hd__a21oi_2 _14217_ (.A1(_04973_),
    .A2(_04976_),
    .B1(_04974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2_2 _14218_ (.A(\b_l[8] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_2 _14219_ (.A(\b_l[7] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05123_));
 sky130_fd_sc_hd__nand2_2 _14220_ (.A(\b_l[6] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05124_));
 sky130_fd_sc_hd__nand2_2 _14221_ (.A(_05123_),
    .B(_05124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_2 _14222_ (.A(\b_l[7] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05126_));
 sky130_fd_sc_hd__and4_2 _14223_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05127_));
 sky130_fd_sc_hd__nand4_2 _14224_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05128_));
 sky130_fd_sc_hd__o221ai_2 _14225_ (.A1(_09264_),
    .A2(_09449_),
    .B1(_05012_),
    .B2(_05126_),
    .C1(_05125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05129_));
 sky130_fd_sc_hd__a21o_2 _14226_ (.A1(_05125_),
    .A2(_05128_),
    .B1(_05122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05130_));
 sky130_fd_sc_hd__a22o_2 _14227_ (.A1(\b_l[8] ),
    .A2(\a_h[7] ),
    .B1(_05125_),
    .B2(_05128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05131_));
 sky130_fd_sc_hd__and4_2 _14228_ (.A(_05125_),
    .B(_05128_),
    .C(\b_l[8] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05132_));
 sky130_fd_sc_hd__o2111ai_2 _14229_ (.A1(_05012_),
    .A2(_05126_),
    .B1(\b_l[8] ),
    .C1(\a_h[7] ),
    .D1(_05125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3b_2 _14230_ (.A_N(_05121_),
    .B(_05129_),
    .C(_05130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_2 _14231_ (.A(_05121_),
    .B(_05131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05135_));
 sky130_fd_sc_hd__nand3_2 _14232_ (.A(_05121_),
    .B(_05131_),
    .C(_05133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05136_));
 sky130_fd_sc_hd__o2bb2ai_2 _14233_ (.A1_N(_05120_),
    .A2_N(_05134_),
    .B1(_05135_),
    .B2(_05132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05137_));
 sky130_fd_sc_hd__a21boi_2 _14234_ (.A1(_05120_),
    .A2(_05134_),
    .B1_N(_05136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05138_));
 sky130_fd_sc_hd__a21oi_2 _14235_ (.A1(_05134_),
    .A2(_05136_),
    .B1(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05139_));
 sky130_fd_sc_hd__a21o_2 _14236_ (.A1(_05134_),
    .A2(_05136_),
    .B1(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05140_));
 sky130_fd_sc_hd__and3_2 _14237_ (.A(_05134_),
    .B(_05136_),
    .C(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05141_));
 sky130_fd_sc_hd__o211ai_2 _14238_ (.A1(_05132_),
    .A2(_05135_),
    .B1(_05134_),
    .C1(_05120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05142_));
 sky130_fd_sc_hd__nand2_2 _14239_ (.A(_05140_),
    .B(_05142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_2 _14240_ (.A(_05139_),
    .B(_05141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05144_));
 sky130_fd_sc_hd__o2bb2ai_2 _14241_ (.A1_N(_04979_),
    .A2_N(_04997_),
    .B1(_04993_),
    .B2(_04990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05145_));
 sky130_fd_sc_hd__a2bb2oi_2 _14242_ (.A1_N(_04990_),
    .A2_N(_04993_),
    .B1(_04997_),
    .B2(_04979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_2 _14243_ (.A(\b_l[5] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_2 _14244_ (.A(\b_l[3] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_2 _14245_ (.A(\b_l[4] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05149_));
 sky130_fd_sc_hd__a22oi_2 _14246_ (.A1(\b_l[4] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_2 _14247_ (.A(_05148_),
    .B(_05149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05151_));
 sky130_fd_sc_hd__nand4_2 _14248_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05152_));
 sky130_fd_sc_hd__a22oi_2 _14249_ (.A1(\b_l[5] ),
    .A2(\a_h[10] ),
    .B1(_05151_),
    .B2(_05152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05153_));
 sky130_fd_sc_hd__o2111a_2 _14250_ (.A1(_02502_),
    .A2(_04182_),
    .B1(\b_l[5] ),
    .C1(\a_h[10] ),
    .D1(_05151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05154_));
 sky130_fd_sc_hd__nor2_2 _14251_ (.A(_05153_),
    .B(_05154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05155_));
 sky130_fd_sc_hd__a21o_2 _14252_ (.A1(_04982_),
    .A2(_04989_),
    .B1(_04985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05156_));
 sky130_fd_sc_hd__a21oi_2 _14253_ (.A1(_04982_),
    .A2(_04989_),
    .B1(_04985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_2 _14254_ (.A(\b_l[2] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_2 _14255_ (.A(\b_l[0] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05159_));
 sky130_fd_sc_hd__a22oi_2 _14256_ (.A1(\b_l[1] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_2 _14257_ (.A(_04988_),
    .B(_05159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_2 _14258_ (.A(\b_l[1] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05162_));
 sky130_fd_sc_hd__nand4_2 _14259_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05163_));
 sky130_fd_sc_hd__o2bb2ai_2 _14260_ (.A1_N(_05161_),
    .A2_N(_05163_),
    .B1(_09155_),
    .B2(_09515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05164_));
 sky130_fd_sc_hd__nand3_2 _14261_ (.A(_05163_),
    .B(\a_h[13] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05165_));
 sky130_fd_sc_hd__nand2_2 _14262_ (.A(_05158_),
    .B(_05163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05166_));
 sky130_fd_sc_hd__a21o_2 _14263_ (.A1(_05161_),
    .A2(_05163_),
    .B1(_05158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05167_));
 sky130_fd_sc_hd__o211ai_2 _14264_ (.A1(_05160_),
    .A2(_05166_),
    .B1(_05156_),
    .C1(_05167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05168_));
 sky130_fd_sc_hd__inv_2 _14265_ (.A(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05169_));
 sky130_fd_sc_hd__o211ai_2 _14266_ (.A1(_05165_),
    .A2(_05160_),
    .B1(_05157_),
    .C1(_05164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05170_));
 sky130_fd_sc_hd__nand2_2 _14267_ (.A(_05168_),
    .B(_05170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05171_));
 sky130_fd_sc_hd__o21ai_2 _14268_ (.A1(_05153_),
    .A2(_05154_),
    .B1(_05171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05172_));
 sky130_fd_sc_hd__nand3_2 _14269_ (.A(_05155_),
    .B(_05168_),
    .C(_05170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05173_));
 sky130_fd_sc_hd__o21ai_2 _14270_ (.A1(_05153_),
    .A2(_05154_),
    .B1(_05170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_2 _14271_ (.A(_05171_),
    .B(_05155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05175_));
 sky130_fd_sc_hd__a21oi_2 _14272_ (.A1(_05172_),
    .A2(_05173_),
    .B1(_05145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05176_));
 sky130_fd_sc_hd__o211ai_2 _14273_ (.A1(_05174_),
    .A2(_05169_),
    .B1(_05146_),
    .C1(_05175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05177_));
 sky130_fd_sc_hd__nand3_2 _14274_ (.A(_05172_),
    .B(_05173_),
    .C(_05145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05178_));
 sky130_fd_sc_hd__nand2_2 _14275_ (.A(_05144_),
    .B(_05177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05179_));
 sky130_fd_sc_hd__o21a_2 _14276_ (.A1(_05139_),
    .A2(_05141_),
    .B1(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05180_));
 sky130_fd_sc_hd__a21oi_2 _14277_ (.A1(_05143_),
    .A2(_05178_),
    .B1(_05176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_2 _14278_ (.A(_05177_),
    .B(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_2 _14279_ (.A1(_05139_),
    .A2(_05141_),
    .B1(_05182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05183_));
 sky130_fd_sc_hd__nand4_2 _14280_ (.A(_05140_),
    .B(_05142_),
    .C(_05177_),
    .D(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05184_));
 sky130_fd_sc_hd__a32oi_2 _14281_ (.A1(_05144_),
    .A2(_05177_),
    .A3(_05178_),
    .B1(_05032_),
    .B2(_05006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05185_));
 sky130_fd_sc_hd__nand3_2 _14282_ (.A(_05033_),
    .B(_05183_),
    .C(_05184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05186_));
 sky130_fd_sc_hd__o211ai_2 _14283_ (.A1(_05139_),
    .A2(_05141_),
    .B1(_05177_),
    .C1(_05178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05187_));
 sky130_fd_sc_hd__a21o_2 _14284_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05188_));
 sky130_fd_sc_hd__a21oi_2 _14285_ (.A1(_05183_),
    .A2(_05184_),
    .B1(_05033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05189_));
 sky130_fd_sc_hd__nand3_2 _14286_ (.A(_05034_),
    .B(_05187_),
    .C(_05188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05190_));
 sky130_fd_sc_hd__and3_2 _14287_ (.A(\a_h[2] ),
    .B(\a_h[3] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05191_));
 sky130_fd_sc_hd__nand4_2 _14288_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[2] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05192_));
 sky130_fd_sc_hd__a22o_2 _14289_ (.A1(\b_l[13] ),
    .A2(\a_h[2] ),
    .B1(\a_h[3] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05193_));
 sky130_fd_sc_hd__and4_2 _14290_ (.A(_05193_),
    .B(\a_h[1] ),
    .C(\b_l[14] ),
    .D(_05192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05194_));
 sky130_fd_sc_hd__o2111ai_2 _14291_ (.A1(_01871_),
    .A2(_05044_),
    .B1(\b_l[14] ),
    .C1(\a_h[1] ),
    .D1(_05193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05195_));
 sky130_fd_sc_hd__a22oi_2 _14292_ (.A1(\b_l[14] ),
    .A2(\a_h[1] ),
    .B1(_05192_),
    .B2(_05193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05196_));
 sky130_fd_sc_hd__a22o_2 _14293_ (.A1(\b_l[14] ),
    .A2(\a_h[1] ),
    .B1(_05192_),
    .B2(_05193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05197_));
 sky130_fd_sc_hd__nor2_2 _14294_ (.A(_05194_),
    .B(_05196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_2 _14295_ (.A(_05195_),
    .B(_05197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05199_));
 sky130_fd_sc_hd__a21oi_2 _14296_ (.A1(_05053_),
    .A2(_05054_),
    .B1(_05052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ai_2 _14297_ (.A1(_04842_),
    .A2(_05056_),
    .B1(_05052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_2 _14298_ (.A(_05055_),
    .B(_05201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05202_));
 sky130_fd_sc_hd__nand2_2 _14299_ (.A(\b_l[11] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05203_));
 sky130_fd_sc_hd__nand2_2 _14300_ (.A(\b_l[9] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05204_));
 sky130_fd_sc_hd__a22oi_2 _14301_ (.A1(\b_l[10] ),
    .A2(\a_h[5] ),
    .B1(\a_h[6] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05205_));
 sky130_fd_sc_hd__nand2_2 _14302_ (.A(_05056_),
    .B(_05204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_2 _14303_ (.A(\b_l[10] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05207_));
 sky130_fd_sc_hd__nand4_2 _14304_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05208_));
 sky130_fd_sc_hd__o2111ai_2 _14305_ (.A1(_05053_),
    .A2(_05207_),
    .B1(\b_l[11] ),
    .C1(\a_h[4] ),
    .D1(_05206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05209_));
 sky130_fd_sc_hd__o2bb2ai_2 _14306_ (.A1_N(_05206_),
    .A2_N(_05208_),
    .B1(_09308_),
    .B2(_09417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05210_));
 sky130_fd_sc_hd__o221ai_2 _14307_ (.A1(_09308_),
    .A2(_09417_),
    .B1(_05053_),
    .B2(_05207_),
    .C1(_05206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05211_));
 sky130_fd_sc_hd__a21o_2 _14308_ (.A1(_05206_),
    .A2(_05208_),
    .B1(_05203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05212_));
 sky130_fd_sc_hd__o211ai_2 _14309_ (.A1(_05057_),
    .A2(_05200_),
    .B1(_05209_),
    .C1(_05210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05213_));
 sky130_fd_sc_hd__a22oi_2 _14310_ (.A1(_05055_),
    .A2(_05201_),
    .B1(_05209_),
    .B2(_05210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05214_));
 sky130_fd_sc_hd__nand3_2 _14311_ (.A(_05212_),
    .B(_05202_),
    .C(_05211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05215_));
 sky130_fd_sc_hd__nand2_2 _14312_ (.A(_05213_),
    .B(_05215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05216_));
 sky130_fd_sc_hd__nand4_2 _14313_ (.A(_05195_),
    .B(_05197_),
    .C(_05213_),
    .D(_05215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05217_));
 sky130_fd_sc_hd__a22o_2 _14314_ (.A1(_05195_),
    .A2(_05197_),
    .B1(_05213_),
    .B2(_05215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05218_));
 sky130_fd_sc_hd__o21ai_2 _14315_ (.A1(_05199_),
    .A2(_05214_),
    .B1(_05213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05219_));
 sky130_fd_sc_hd__o21a_2 _14316_ (.A1(_05199_),
    .A2(_05214_),
    .B1(_05213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05220_));
 sky130_fd_sc_hd__o211ai_2 _14317_ (.A1(_05194_),
    .A2(_05196_),
    .B1(_05213_),
    .C1(_05215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_2 _14318_ (.A(_05216_),
    .B(_05198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05222_));
 sky130_fd_sc_hd__nand3_2 _14319_ (.A(_05024_),
    .B(_05221_),
    .C(_05222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05223_));
 sky130_fd_sc_hd__nand3_2 _14320_ (.A(_05218_),
    .B(_05023_),
    .C(_05217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_2 _14321_ (.A(_05223_),
    .B(_05224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05225_));
 sky130_fd_sc_hd__o21a_2 _14322_ (.A1(_05050_),
    .A2(_05065_),
    .B1(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05226_));
 sky130_fd_sc_hd__o21ai_2 _14323_ (.A1(_05050_),
    .A2(_05065_),
    .B1(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05227_));
 sky130_fd_sc_hd__and3_2 _14324_ (.A(_05223_),
    .B(_05224_),
    .C(_05227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05228_));
 sky130_fd_sc_hd__nand3_2 _14325_ (.A(_05223_),
    .B(_05224_),
    .C(_05227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05229_));
 sky130_fd_sc_hd__o211a_2 _14326_ (.A1(_05050_),
    .A2(_05065_),
    .B1(_05225_),
    .C1(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05230_));
 sky130_fd_sc_hd__nand2_2 _14327_ (.A(_05225_),
    .B(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05231_));
 sky130_fd_sc_hd__a21oi_2 _14328_ (.A1(_05223_),
    .A2(_05224_),
    .B1(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05232_));
 sky130_fd_sc_hd__a21o_2 _14329_ (.A1(_05223_),
    .A2(_05224_),
    .B1(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05233_));
 sky130_fd_sc_hd__and3_2 _14330_ (.A(_05223_),
    .B(_05224_),
    .C(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05234_));
 sky130_fd_sc_hd__o2111ai_2 _14331_ (.A1(_05050_),
    .A2(_05065_),
    .B1(_05223_),
    .C1(_05224_),
    .D1(_05063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_2 _14332_ (.A(_05233_),
    .B(_05235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_2 _14333_ (.A(_05229_),
    .B(_05231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05237_));
 sky130_fd_sc_hd__o211ai_2 _14334_ (.A1(_05232_),
    .A2(_05234_),
    .B1(_05186_),
    .C1(_05190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05238_));
 sky130_fd_sc_hd__inv_2 _14335_ (.A(_05238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05239_));
 sky130_fd_sc_hd__o2bb2ai_2 _14336_ (.A1_N(_05186_),
    .A2_N(_05190_),
    .B1(_05228_),
    .B2(_05230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_2 _14337_ (.A(_05119_),
    .B(_05240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05241_));
 sky130_fd_sc_hd__nand3_2 _14338_ (.A(_05119_),
    .B(_05238_),
    .C(_05240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05242_));
 sky130_fd_sc_hd__nand4_2 _14339_ (.A(_05186_),
    .B(_05190_),
    .C(_05233_),
    .D(_05235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05243_));
 sky130_fd_sc_hd__o2bb2ai_2 _14340_ (.A1_N(_05186_),
    .A2_N(_05190_),
    .B1(_05232_),
    .B2(_05234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05244_));
 sky130_fd_sc_hd__nand3_2 _14341_ (.A(_05244_),
    .B(_05118_),
    .C(_05243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_2 _14342_ (.A(_05242_),
    .B(_05245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05246_));
 sky130_fd_sc_hd__o211ai_2 _14343_ (.A1(_05239_),
    .A2(_05241_),
    .B1(_05245_),
    .C1(_05116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05247_));
 sky130_fd_sc_hd__a21o_2 _14344_ (.A1(_05242_),
    .A2(_05245_),
    .B1(_05116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05248_));
 sky130_fd_sc_hd__nand3_2 _14345_ (.A(_05107_),
    .B(_05247_),
    .C(_05248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05249_));
 sky130_fd_sc_hd__nand3b_2 _14346_ (.A_N(_05116_),
    .B(_05242_),
    .C(_05245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_2 _14347_ (.A(_05246_),
    .B(_05116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05251_));
 sky130_fd_sc_hd__nand3_2 _14348_ (.A(_05251_),
    .B(_05106_),
    .C(_05250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05252_));
 sky130_fd_sc_hd__nand3_2 _14349_ (.A(_05249_),
    .B(_05252_),
    .C(_05088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05253_));
 sky130_fd_sc_hd__o2bb2ai_2 _14350_ (.A1_N(_05249_),
    .A2_N(_05252_),
    .B1(_04837_),
    .B2(_05087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05254_));
 sky130_fd_sc_hd__a21oi_2 _14351_ (.A1(_05253_),
    .A2(_05254_),
    .B1(_05096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05255_));
 sky130_fd_sc_hd__nand3_2 _14352_ (.A(_05254_),
    .B(_05096_),
    .C(_05253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2b_2 _14353_ (.A_N(_05255_),
    .B(_05256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05257_));
 sky130_fd_sc_hd__a21oi_2 _14354_ (.A1(_05100_),
    .A2(_05105_),
    .B1(_05257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05258_));
 sky130_fd_sc_hd__a31o_2 _14355_ (.A1(_05100_),
    .A2(_05105_),
    .A3(_05257_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05259_));
 sky130_fd_sc_hd__nor2_2 _14356_ (.A(_05258_),
    .B(_05259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00321_));
 sky130_fd_sc_hd__o21ai_2 _14357_ (.A1(_05098_),
    .A2(_05255_),
    .B1(_05256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05260_));
 sky130_fd_sc_hd__and2_2 _14358_ (.A(_05100_),
    .B(_05256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05261_));
 sky130_fd_sc_hd__o211ai_2 _14359_ (.A1(_04831_),
    .A2(_05102_),
    .B1(_05261_),
    .C1(_05101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_2 _14360_ (.A(_05262_),
    .B(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05263_));
 sky130_fd_sc_hd__a32oi_2 _14361_ (.A1(_05107_),
    .A2(_05247_),
    .A3(_05248_),
    .B1(_05252_),
    .B2(_05089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05264_));
 sky130_fd_sc_hd__and3_2 _14362_ (.A(_05112_),
    .B(\b_l[15] ),
    .C(\a_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05265_));
 sky130_fd_sc_hd__a32oi_2 _14363_ (.A1(_05119_),
    .A2(_05238_),
    .A3(_05240_),
    .B1(_05245_),
    .B2(_05116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05266_));
 sky130_fd_sc_hd__o2bb2ai_2 _14364_ (.A1_N(_05116_),
    .A2_N(_05245_),
    .B1(_05239_),
    .B2(_05241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05267_));
 sky130_fd_sc_hd__a22oi_2 _14365_ (.A1(_05183_),
    .A2(_05185_),
    .B1(_05190_),
    .B2(_05237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05268_));
 sky130_fd_sc_hd__a21oi_2 _14366_ (.A1(_05186_),
    .A2(_05236_),
    .B1(_05189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2_2 _14367_ (.A(\b_l[5] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_2 _14368_ (.A(\b_l[3] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_2 _14369_ (.A(\b_l[4] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05272_));
 sky130_fd_sc_hd__a22oi_2 _14370_ (.A1(\b_l[4] ),
    .A2(\a_h[12] ),
    .B1(\a_h[13] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05273_));
 sky130_fd_sc_hd__nand2_2 _14371_ (.A(_05271_),
    .B(_05272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05274_));
 sky130_fd_sc_hd__nand4_2 _14372_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05275_));
 sky130_fd_sc_hd__o221a_2 _14373_ (.A1(_09220_),
    .A2(_09493_),
    .B1(_02613_),
    .B2(_04182_),
    .C1(_05274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05276_));
 sky130_fd_sc_hd__o221ai_2 _14374_ (.A1(_09220_),
    .A2(_09493_),
    .B1(_02613_),
    .B2(_04182_),
    .C1(_05274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05277_));
 sky130_fd_sc_hd__a21oi_2 _14375_ (.A1(_05274_),
    .A2(_05275_),
    .B1(_05270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05278_));
 sky130_fd_sc_hd__a21o_2 _14376_ (.A1(_05274_),
    .A2(_05275_),
    .B1(_05270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05279_));
 sky130_fd_sc_hd__a22o_2 _14377_ (.A1(\b_l[5] ),
    .A2(\a_h[11] ),
    .B1(_05274_),
    .B2(_05275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05280_));
 sky130_fd_sc_hd__o2111ai_2 _14378_ (.A1(_02613_),
    .A2(_04182_),
    .B1(\b_l[5] ),
    .C1(\a_h[11] ),
    .D1(_05274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05281_));
 sky130_fd_sc_hd__nand2_2 _14379_ (.A(_05280_),
    .B(_05281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05282_));
 sky130_fd_sc_hd__nand2_2 _14380_ (.A(\b_l[2] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05283_));
 sky130_fd_sc_hd__nand2_2 _14381_ (.A(_05162_),
    .B(_05283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2_2 _14382_ (.A(\b_l[2] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05285_));
 sky130_fd_sc_hd__nand4_2 _14383_ (.A(\b_l[1] ),
    .B(\b_l[2] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05286_));
 sky130_fd_sc_hd__o21ai_2 _14384_ (.A1(_04988_),
    .A2(_05285_),
    .B1(_05284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05287_));
 sky130_fd_sc_hd__o211ai_2 _14385_ (.A1(_05158_),
    .A2(_05160_),
    .B1(_05163_),
    .C1(_05287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05288_));
 sky130_fd_sc_hd__nand4_2 _14386_ (.A(_05161_),
    .B(_05166_),
    .C(_05284_),
    .D(_05286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_2 _14387_ (.A(_05288_),
    .B(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_2 _14388_ (.A(_05277_),
    .B(_05279_),
    .C(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05291_));
 sky130_fd_sc_hd__nand4_2 _14389_ (.A(_05277_),
    .B(_05279_),
    .C(_05288_),
    .D(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05292_));
 sky130_fd_sc_hd__o21ai_2 _14390_ (.A1(_05276_),
    .A2(_05278_),
    .B1(_05290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05293_));
 sky130_fd_sc_hd__nand4_2 _14391_ (.A(_05280_),
    .B(_05281_),
    .C(_05288_),
    .D(_05289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05294_));
 sky130_fd_sc_hd__nand2_2 _14392_ (.A(_05290_),
    .B(_05282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_2 _14393_ (.A(_05155_),
    .B(_05168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05296_));
 sky130_fd_sc_hd__nand4_2 _14394_ (.A(_05170_),
    .B(_05292_),
    .C(_05293_),
    .D(_05296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05297_));
 sky130_fd_sc_hd__nand4_2 _14395_ (.A(_05168_),
    .B(_05174_),
    .C(_05294_),
    .D(_05295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05298_));
 sky130_fd_sc_hd__a21o_2 _14396_ (.A1(_05147_),
    .A2(_05152_),
    .B1(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05299_));
 sky130_fd_sc_hd__a21oi_2 _14397_ (.A1(_05147_),
    .A2(_05152_),
    .B1(_05150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_2 _14398_ (.A(\b_l[8] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05301_));
 sky130_fd_sc_hd__nand2_2 _14399_ (.A(\b_l[6] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05302_));
 sky130_fd_sc_hd__nand2_2 _14400_ (.A(_05126_),
    .B(_05302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05303_));
 sky130_fd_sc_hd__nand3_2 _14401_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05304_));
 sky130_fd_sc_hd__and3_2 _14402_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(_04259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05305_));
 sky130_fd_sc_hd__nand4_2 _14403_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05306_));
 sky130_fd_sc_hd__a21oi_2 _14404_ (.A1(_05303_),
    .A2(_05306_),
    .B1(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05307_));
 sky130_fd_sc_hd__a21o_2 _14405_ (.A1(_05303_),
    .A2(_05306_),
    .B1(_05301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05308_));
 sky130_fd_sc_hd__o221a_2 _14406_ (.A1(_09264_),
    .A2(_09460_),
    .B1(_09482_),
    .B2(_05304_),
    .C1(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05309_));
 sky130_fd_sc_hd__o221ai_2 _14407_ (.A1(_09264_),
    .A2(_09460_),
    .B1(_09482_),
    .B2(_05304_),
    .C1(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05310_));
 sky130_fd_sc_hd__a21oi_2 _14408_ (.A1(_05308_),
    .A2(_05310_),
    .B1(_05299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_2 _14409_ (.A1(_05307_),
    .A2(_05309_),
    .B1(_05300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05312_));
 sky130_fd_sc_hd__nand3_2 _14410_ (.A(_05308_),
    .B(_05310_),
    .C(_05299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05313_));
 sky130_fd_sc_hd__a31o_2 _14411_ (.A1(\b_l[8] ),
    .A2(_05125_),
    .A3(\a_h[7] ),
    .B1(_05127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05314_));
 sky130_fd_sc_hd__o31a_2 _14412_ (.A1(_09460_),
    .A2(_09471_),
    .A3(_04260_),
    .B1(_05133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05315_));
 sky130_fd_sc_hd__a21oi_2 _14413_ (.A1(_05312_),
    .A2(_05313_),
    .B1(_05315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05316_));
 sky130_fd_sc_hd__and3_2 _14414_ (.A(_05312_),
    .B(_05313_),
    .C(_05315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05317_));
 sky130_fd_sc_hd__a21oi_2 _14415_ (.A1(_05312_),
    .A2(_05313_),
    .B1(_05314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05318_));
 sky130_fd_sc_hd__o21ai_2 _14416_ (.A1(_05127_),
    .A2(_05132_),
    .B1(_05313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05319_));
 sky130_fd_sc_hd__o311a_2 _14417_ (.A1(_05300_),
    .A2(_05307_),
    .A3(_05309_),
    .B1(_05314_),
    .C1(_05312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05320_));
 sky130_fd_sc_hd__o2bb2ai_2 _14418_ (.A1_N(_05297_),
    .A2_N(_05298_),
    .B1(_05318_),
    .B2(_05320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05321_));
 sky130_fd_sc_hd__o21ai_2 _14419_ (.A1(_05316_),
    .A2(_05317_),
    .B1(_05297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05322_));
 sky130_fd_sc_hd__o211ai_2 _14420_ (.A1(_05316_),
    .A2(_05317_),
    .B1(_05297_),
    .C1(_05298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05323_));
 sky130_fd_sc_hd__nand3_2 _14421_ (.A(_05177_),
    .B(_05321_),
    .C(_05323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05324_));
 sky130_fd_sc_hd__nand3_2 _14422_ (.A(_05181_),
    .B(_05321_),
    .C(_05323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05325_));
 sky130_fd_sc_hd__o211ai_2 _14423_ (.A1(_05318_),
    .A2(_05320_),
    .B1(_05297_),
    .C1(_05298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05326_));
 sky130_fd_sc_hd__o2bb2ai_2 _14424_ (.A1_N(_05297_),
    .A2_N(_05298_),
    .B1(_05316_),
    .B2(_05317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05327_));
 sky130_fd_sc_hd__a21oi_2 _14425_ (.A1(_05321_),
    .A2(_05323_),
    .B1(_05181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05328_));
 sky130_fd_sc_hd__nand4_2 _14426_ (.A(_05178_),
    .B(_05179_),
    .C(_05326_),
    .D(_05327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05329_));
 sky130_fd_sc_hd__nand2_2 _14427_ (.A(\b_l[12] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_2 _14428_ (.A(\b_l[13] ),
    .B(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05331_));
 sky130_fd_sc_hd__nand2_2 _14429_ (.A(_05330_),
    .B(_05331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05332_));
 sky130_fd_sc_hd__nand2_2 _14430_ (.A(\b_l[13] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05333_));
 sky130_fd_sc_hd__nand4_2 _14431_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[3] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05334_));
 sky130_fd_sc_hd__and2_2 _14432_ (.A(\b_l[14] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05335_));
 sky130_fd_sc_hd__and3_2 _14433_ (.A(_05332_),
    .B(_05335_),
    .C(_05334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05336_));
 sky130_fd_sc_hd__o2111ai_2 _14434_ (.A1(_01888_),
    .A2(_05044_),
    .B1(\b_l[14] ),
    .C1(\a_h[2] ),
    .D1(_05332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05337_));
 sky130_fd_sc_hd__a21oi_2 _14435_ (.A1(_05332_),
    .A2(_05334_),
    .B1(_05335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05338_));
 sky130_fd_sc_hd__a22o_2 _14436_ (.A1(\b_l[14] ),
    .A2(\a_h[2] ),
    .B1(_05332_),
    .B2(_05334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05339_));
 sky130_fd_sc_hd__nor2_2 _14437_ (.A(_05336_),
    .B(_05338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05340_));
 sky130_fd_sc_hd__a21o_2 _14438_ (.A1(_05203_),
    .A2(_05208_),
    .B1(_05205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05341_));
 sky130_fd_sc_hd__a21oi_2 _14439_ (.A1(_05203_),
    .A2(_05208_),
    .B1(_05205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05342_));
 sky130_fd_sc_hd__nand2_2 _14440_ (.A(\b_l[11] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05343_));
 sky130_fd_sc_hd__nand2_2 _14441_ (.A(\b_l[9] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05344_));
 sky130_fd_sc_hd__a22oi_2 _14442_ (.A1(\b_l[10] ),
    .A2(\a_h[6] ),
    .B1(\a_h[7] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_2 _14443_ (.A(_05207_),
    .B(_05344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05346_));
 sky130_fd_sc_hd__nand2_2 _14444_ (.A(\b_l[10] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05347_));
 sky130_fd_sc_hd__nand4_2 _14445_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[6] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05348_));
 sky130_fd_sc_hd__nand3_2 _14446_ (.A(_05348_),
    .B(\a_h[5] ),
    .C(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05349_));
 sky130_fd_sc_hd__o2bb2ai_2 _14447_ (.A1_N(_05346_),
    .A2_N(_05348_),
    .B1(_09308_),
    .B2(_09428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05350_));
 sky130_fd_sc_hd__a21o_2 _14448_ (.A1(_05346_),
    .A2(_05348_),
    .B1(_05343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05351_));
 sky130_fd_sc_hd__o221ai_2 _14449_ (.A1(_09308_),
    .A2(_09428_),
    .B1(_05204_),
    .B2(_05347_),
    .C1(_05346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05352_));
 sky130_fd_sc_hd__o211ai_2 _14450_ (.A1(_05349_),
    .A2(_05345_),
    .B1(_05342_),
    .C1(_05350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05353_));
 sky130_fd_sc_hd__nand3_2 _14451_ (.A(_05351_),
    .B(_05352_),
    .C(_05341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_2 _14452_ (.A(_05353_),
    .B(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_2 _14453_ (.A(_05355_),
    .B(_05340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05356_));
 sky130_fd_sc_hd__o211ai_2 _14454_ (.A1(_05336_),
    .A2(_05338_),
    .B1(_05353_),
    .C1(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05357_));
 sky130_fd_sc_hd__nand2_2 _14455_ (.A(_05340_),
    .B(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05358_));
 sky130_fd_sc_hd__nand4_2 _14456_ (.A(_05337_),
    .B(_05339_),
    .C(_05353_),
    .D(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05359_));
 sky130_fd_sc_hd__a22o_2 _14457_ (.A1(_05337_),
    .A2(_05339_),
    .B1(_05353_),
    .B2(_05354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05360_));
 sky130_fd_sc_hd__and3_2 _14458_ (.A(_05360_),
    .B(_05137_),
    .C(_05359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05361_));
 sky130_fd_sc_hd__nand3_2 _14459_ (.A(_05360_),
    .B(_05137_),
    .C(_05359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05362_));
 sky130_fd_sc_hd__nand3_2 _14460_ (.A(_05138_),
    .B(_05356_),
    .C(_05357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05363_));
 sky130_fd_sc_hd__a21oi_2 _14461_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05364_));
 sky130_fd_sc_hd__and3_2 _14462_ (.A(_05220_),
    .B(_05362_),
    .C(_05363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05365_));
 sky130_fd_sc_hd__a21oi_2 _14463_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05366_));
 sky130_fd_sc_hd__a21o_2 _14464_ (.A1(_05362_),
    .A2(_05363_),
    .B1(_05219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05367_));
 sky130_fd_sc_hd__a31oi_2 _14465_ (.A1(_05138_),
    .A2(_05356_),
    .A3(_05357_),
    .B1(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05368_));
 sky130_fd_sc_hd__a31o_2 _14466_ (.A1(_05138_),
    .A2(_05356_),
    .A3(_05357_),
    .B1(_05220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05369_));
 sky130_fd_sc_hd__and3_2 _14467_ (.A(_05362_),
    .B(_05363_),
    .C(_05219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05370_));
 sky130_fd_sc_hd__o21ai_2 _14468_ (.A1(_05361_),
    .A2(_05369_),
    .B1(_05367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05371_));
 sky130_fd_sc_hd__a21oi_2 _14469_ (.A1(_05362_),
    .A2(_05368_),
    .B1(_05366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05372_));
 sky130_fd_sc_hd__o221ai_2 _14470_ (.A1(_05366_),
    .A2(_05370_),
    .B1(_05180_),
    .B2(_05324_),
    .C1(_05329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05373_));
 sky130_fd_sc_hd__o2bb2ai_2 _14471_ (.A1_N(_05325_),
    .A2_N(_05329_),
    .B1(_05364_),
    .B2(_05365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05374_));
 sky130_fd_sc_hd__o2bb2ai_2 _14472_ (.A1_N(_05325_),
    .A2_N(_05329_),
    .B1(_05366_),
    .B2(_05370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05375_));
 sky130_fd_sc_hd__o211ai_2 _14473_ (.A1(_05364_),
    .A2(_05365_),
    .B1(_05325_),
    .C1(_05329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05376_));
 sky130_fd_sc_hd__nand3_2 _14474_ (.A(_05268_),
    .B(_05373_),
    .C(_05374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05377_));
 sky130_fd_sc_hd__nand3_2 _14475_ (.A(_05269_),
    .B(_05375_),
    .C(_05376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_2 _14476_ (.A(\b_l[15] ),
    .B(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05379_));
 sky130_fd_sc_hd__a31o_2 _14477_ (.A1(\b_l[14] ),
    .A2(\a_h[1] ),
    .A3(_05193_),
    .B1(_05191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05380_));
 sky130_fd_sc_hd__a31o_2 _14478_ (.A1(_05217_),
    .A2(_05218_),
    .A3(_05023_),
    .B1(_05226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05381_));
 sky130_fd_sc_hd__a31o_2 _14479_ (.A1(_05024_),
    .A2(_05221_),
    .A3(_05222_),
    .B1(_05227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05382_));
 sky130_fd_sc_hd__o211ai_2 _14480_ (.A1(_05191_),
    .A2(_05194_),
    .B1(_05223_),
    .C1(_05381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05383_));
 sky130_fd_sc_hd__inv_2 _14481_ (.A(_05383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05384_));
 sky130_fd_sc_hd__o2111ai_2 _14482_ (.A1(_01871_),
    .A2(_05044_),
    .B1(_05195_),
    .C1(_05224_),
    .D1(_05382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05385_));
 sky130_fd_sc_hd__a31oi_2 _14483_ (.A1(_05223_),
    .A2(_05380_),
    .A3(_05381_),
    .B1(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05386_));
 sky130_fd_sc_hd__and4_2 _14484_ (.A(_05383_),
    .B(_05385_),
    .C(\b_l[15] ),
    .D(\a_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05387_));
 sky130_fd_sc_hd__a22oi_2 _14485_ (.A1(\b_l[15] ),
    .A2(\a_h[1] ),
    .B1(_05383_),
    .B2(_05385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05388_));
 sky130_fd_sc_hd__and3_2 _14486_ (.A(_05379_),
    .B(_05383_),
    .C(_05385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05389_));
 sky130_fd_sc_hd__a21oi_2 _14487_ (.A1(_05383_),
    .A2(_05385_),
    .B1(_05379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05390_));
 sky130_fd_sc_hd__a21oi_2 _14488_ (.A1(_05385_),
    .A2(_05386_),
    .B1(_05388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05391_));
 sky130_fd_sc_hd__o2bb2ai_2 _14489_ (.A1_N(_05377_),
    .A2_N(_05378_),
    .B1(_05389_),
    .B2(_05390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05392_));
 sky130_fd_sc_hd__o211ai_2 _14490_ (.A1(_05387_),
    .A2(_05388_),
    .B1(_05377_),
    .C1(_05378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05393_));
 sky130_fd_sc_hd__nand3_2 _14491_ (.A(_05267_),
    .B(_05392_),
    .C(_05393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05394_));
 sky130_fd_sc_hd__inv_2 _14492_ (.A(_05394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_2 _14493_ (.A(_05377_),
    .B(_05391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05396_));
 sky130_fd_sc_hd__o211ai_2 _14494_ (.A1(_05389_),
    .A2(_05390_),
    .B1(_05377_),
    .C1(_05378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05397_));
 sky130_fd_sc_hd__o2bb2ai_2 _14495_ (.A1_N(_05377_),
    .A2_N(_05378_),
    .B1(_05387_),
    .B2(_05388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05398_));
 sky130_fd_sc_hd__nand3_2 _14496_ (.A(_05266_),
    .B(_05397_),
    .C(_05398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05399_));
 sky130_fd_sc_hd__o21ai_2 _14497_ (.A1(_05110_),
    .A2(_05265_),
    .B1(_05394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05400_));
 sky130_fd_sc_hd__o211a_2 _14498_ (.A1(_05110_),
    .A2(_05265_),
    .B1(_05394_),
    .C1(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05401_));
 sky130_fd_sc_hd__o211ai_2 _14499_ (.A1(_05110_),
    .A2(_05265_),
    .B1(_05394_),
    .C1(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05402_));
 sky130_fd_sc_hd__a2bb2oi_2 _14500_ (.A1_N(_05111_),
    .A2_N(_05113_),
    .B1(_05394_),
    .B2(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05403_));
 sky130_fd_sc_hd__o21a_2 _14501_ (.A1(_05111_),
    .A2(_05113_),
    .B1(_05399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_2 _14502_ (.A(_05399_),
    .B(_05400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05405_));
 sky130_fd_sc_hd__o21ba_2 _14503_ (.A1(_05401_),
    .A2(_05403_),
    .B1_N(_05264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05406_));
 sky130_fd_sc_hd__o21bai_2 _14504_ (.A1(_05401_),
    .A2(_05403_),
    .B1_N(_05264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05407_));
 sky130_fd_sc_hd__nand3b_2 _14505_ (.A_N(_05403_),
    .B(_05264_),
    .C(_05402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_2 _14506_ (.A(_05407_),
    .B(_05408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05409_));
 sky130_fd_sc_hd__a21oi_2 _14507_ (.A1(_05263_),
    .A2(_05409_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05410_));
 sky130_fd_sc_hd__o21a_2 _14508_ (.A1(_05263_),
    .A2(_05409_),
    .B1(_05410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00322_));
 sky130_fd_sc_hd__a32oi_2 _14509_ (.A1(_05269_),
    .A2(_05375_),
    .A3(_05376_),
    .B1(_05377_),
    .B2(_05391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_2 _14510_ (.A(_05378_),
    .B(_05396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05412_));
 sky130_fd_sc_hd__a2bb2oi_2 _14511_ (.A1_N(_05180_),
    .A2_N(_05324_),
    .B1(_05329_),
    .B2(_05372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05413_));
 sky130_fd_sc_hd__o22ai_2 _14512_ (.A1(_05324_),
    .A2(_05180_),
    .B1(_05371_),
    .B2(_05328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05414_));
 sky130_fd_sc_hd__o21ai_2 _14513_ (.A1(_05318_),
    .A2(_05320_),
    .B1(_05298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05415_));
 sky130_fd_sc_hd__o21ai_2 _14514_ (.A1(_05270_),
    .A2(_05273_),
    .B1(_05275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05416_));
 sky130_fd_sc_hd__o22a_2 _14515_ (.A1(_02613_),
    .A2(_04182_),
    .B1(_05270_),
    .B2(_05273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05417_));
 sky130_fd_sc_hd__nand2_2 _14516_ (.A(\b_l[8] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05418_));
 sky130_fd_sc_hd__nand2_2 _14517_ (.A(\b_l[7] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_2 _14518_ (.A(\b_l[6] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_2 _14519_ (.A(_05419_),
    .B(_05420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05421_));
 sky130_fd_sc_hd__nand4_2 _14520_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05422_));
 sky130_fd_sc_hd__a21o_2 _14521_ (.A1(_05421_),
    .A2(_05422_),
    .B1(_05418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05423_));
 sky130_fd_sc_hd__o311a_2 _14522_ (.A1(_09482_),
    .A2(_09493_),
    .A3(_04260_),
    .B1(_05418_),
    .C1(_05421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05424_));
 sky130_fd_sc_hd__o211ai_2 _14523_ (.A1(_09264_),
    .A2(_09471_),
    .B1(_05421_),
    .C1(_05422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05425_));
 sky130_fd_sc_hd__nand4_2 _14524_ (.A(_05421_),
    .B(_05422_),
    .C(\b_l[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05426_));
 sky130_fd_sc_hd__a22o_2 _14525_ (.A1(\b_l[8] ),
    .A2(\a_h[9] ),
    .B1(_05421_),
    .B2(_05422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05427_));
 sky130_fd_sc_hd__nand3_2 _14526_ (.A(_05427_),
    .B(_05416_),
    .C(_05426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05428_));
 sky130_fd_sc_hd__nand2_2 _14527_ (.A(_05417_),
    .B(_05423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05429_));
 sky130_fd_sc_hd__nand3_2 _14528_ (.A(_05417_),
    .B(_05423_),
    .C(_05425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05430_));
 sky130_fd_sc_hd__and3_2 _14529_ (.A(_05303_),
    .B(\a_h[8] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05431_));
 sky130_fd_sc_hd__a21bo_2 _14530_ (.A1(_05301_),
    .A2(_05306_),
    .B1_N(_05303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05432_));
 sky130_fd_sc_hd__o211ai_2 _14531_ (.A1(_05424_),
    .A2(_05429_),
    .B1(_05432_),
    .C1(_05428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05433_));
 sky130_fd_sc_hd__o2bb2ai_2 _14532_ (.A1_N(_05428_),
    .A2_N(_05430_),
    .B1(_05431_),
    .B2(_05305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05434_));
 sky130_fd_sc_hd__a21boi_2 _14533_ (.A1(_05428_),
    .A2(_05430_),
    .B1_N(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05435_));
 sky130_fd_sc_hd__o211a_2 _14534_ (.A1(_05305_),
    .A2(_05431_),
    .B1(_05430_),
    .C1(_05428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05436_));
 sky130_fd_sc_hd__nand2_2 _14535_ (.A(_05433_),
    .B(_05434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05437_));
 sky130_fd_sc_hd__nand3_2 _14536_ (.A(_05280_),
    .B(_05281_),
    .C(_05288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05438_));
 sky130_fd_sc_hd__and3_2 _14537_ (.A(_04988_),
    .B(\a_h[15] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05439_));
 sky130_fd_sc_hd__nor2_2 _14538_ (.A(_09220_),
    .B(_09504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_2 _14539_ (.A(\b_l[5] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05441_));
 sky130_fd_sc_hd__nand2_2 _14540_ (.A(\b_l[3] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_2 _14541_ (.A(\b_l[4] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05443_));
 sky130_fd_sc_hd__a22oi_2 _14542_ (.A1(\b_l[4] ),
    .A2(\a_h[13] ),
    .B1(\a_h[14] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05444_));
 sky130_fd_sc_hd__nand2_2 _14543_ (.A(_05442_),
    .B(_05443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05445_));
 sky130_fd_sc_hd__nand2_2 _14544_ (.A(\b_l[4] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05446_));
 sky130_fd_sc_hd__o2bb2ai_2 _14545_ (.A1_N(_05442_),
    .A2_N(_05443_),
    .B1(_05446_),
    .B2(_05271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05447_));
 sky130_fd_sc_hd__o221ai_2 _14546_ (.A1(_09220_),
    .A2(_09504_),
    .B1(_05271_),
    .B2(_05446_),
    .C1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05448_));
 sky130_fd_sc_hd__nand2_2 _14547_ (.A(_05447_),
    .B(_05440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05449_));
 sky130_fd_sc_hd__o2111ai_2 _14548_ (.A1(_05271_),
    .A2(_05446_),
    .B1(\b_l[5] ),
    .C1(\a_h[12] ),
    .D1(_05445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_2 _14549_ (.A1(_09220_),
    .A2(_09504_),
    .B1(_05447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05451_));
 sky130_fd_sc_hd__nand3_2 _14550_ (.A(_05451_),
    .B(_05439_),
    .C(_05450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05452_));
 sky130_fd_sc_hd__o211ai_2 _14551_ (.A1(_04987_),
    .A2(_05285_),
    .B1(_05448_),
    .C1(_05449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_2 _14552_ (.A(_05452_),
    .B(_05453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05454_));
 sky130_fd_sc_hd__a21oi_2 _14553_ (.A1(_05289_),
    .A2(_05438_),
    .B1(_05454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05455_));
 sky130_fd_sc_hd__nand4_2 _14554_ (.A(_05288_),
    .B(_05291_),
    .C(_05452_),
    .D(_05453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05456_));
 sky130_fd_sc_hd__a22oi_2 _14555_ (.A1(_05288_),
    .A2(_05291_),
    .B1(_05452_),
    .B2(_05453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05457_));
 sky130_fd_sc_hd__nand3_2 _14556_ (.A(_05289_),
    .B(_05438_),
    .C(_05454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05458_));
 sky130_fd_sc_hd__nand3_2 _14557_ (.A(_05437_),
    .B(_05456_),
    .C(_05458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05459_));
 sky130_fd_sc_hd__o22ai_2 _14558_ (.A1(_05435_),
    .A2(_05436_),
    .B1(_05455_),
    .B2(_05457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05460_));
 sky130_fd_sc_hd__nand4_2 _14559_ (.A(_05433_),
    .B(_05434_),
    .C(_05456_),
    .D(_05458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05461_));
 sky130_fd_sc_hd__o21ai_2 _14560_ (.A1(_05455_),
    .A2(_05457_),
    .B1(_05437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05462_));
 sky130_fd_sc_hd__nand4_2 _14561_ (.A(_05298_),
    .B(_05322_),
    .C(_05461_),
    .D(_05462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05463_));
 sky130_fd_sc_hd__nand4_2 _14562_ (.A(_05297_),
    .B(_05415_),
    .C(_05459_),
    .D(_05460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05464_));
 sky130_fd_sc_hd__nand2_2 _14563_ (.A(_05463_),
    .B(_05464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05465_));
 sky130_fd_sc_hd__nand2_2 _14564_ (.A(\b_l[13] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05466_));
 sky130_fd_sc_hd__nand2_2 _14565_ (.A(\b_l[12] ),
    .B(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05467_));
 sky130_fd_sc_hd__and4_2 _14566_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05468_));
 sky130_fd_sc_hd__nand4_2 _14567_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[4] ),
    .D(\a_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_2 _14568_ (.A(_05333_),
    .B(_05467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05470_));
 sky130_fd_sc_hd__and4_2 _14569_ (.A(_05470_),
    .B(\a_h[3] ),
    .C(\b_l[14] ),
    .D(_05469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05471_));
 sky130_fd_sc_hd__o2111ai_2 _14570_ (.A1(_05330_),
    .A2(_05466_),
    .B1(\b_l[14] ),
    .C1(\a_h[3] ),
    .D1(_05470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05472_));
 sky130_fd_sc_hd__o2bb2a_2 _14571_ (.A1_N(_05469_),
    .A2_N(_05470_),
    .B1(_09362_),
    .B2(_09406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05473_));
 sky130_fd_sc_hd__a22o_2 _14572_ (.A1(\b_l[14] ),
    .A2(\a_h[3] ),
    .B1(_05469_),
    .B2(_05470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05474_));
 sky130_fd_sc_hd__nor2_2 _14573_ (.A(_05471_),
    .B(_05473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_2 _14574_ (.A(_05472_),
    .B(_05474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05476_));
 sky130_fd_sc_hd__a21oi_2 _14575_ (.A1(_05343_),
    .A2(_05348_),
    .B1(_05345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_2 _14576_ (.A(\b_l[11] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_2 _14577_ (.A(\b_l[9] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_2 _14578_ (.A(_05347_),
    .B(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05480_));
 sky130_fd_sc_hd__nand4_2 _14579_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05481_));
 sky130_fd_sc_hd__a21o_2 _14580_ (.A1(_05480_),
    .A2(_05481_),
    .B1(_05478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05482_));
 sky130_fd_sc_hd__o211ai_2 _14581_ (.A1(_09308_),
    .A2(_09439_),
    .B1(_05480_),
    .C1(_05481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05483_));
 sky130_fd_sc_hd__o2bb2ai_2 _14582_ (.A1_N(_05480_),
    .A2_N(_05481_),
    .B1(_09308_),
    .B2(_09439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05484_));
 sky130_fd_sc_hd__nand4_2 _14583_ (.A(_05480_),
    .B(_05481_),
    .C(\b_l[11] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05485_));
 sky130_fd_sc_hd__nand3b_2 _14584_ (.A_N(_05477_),
    .B(_05482_),
    .C(_05483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05486_));
 sky130_fd_sc_hd__nand3_2 _14585_ (.A(_05477_),
    .B(_05484_),
    .C(_05485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05487_));
 sky130_fd_sc_hd__a22o_2 _14586_ (.A1(_05472_),
    .A2(_05474_),
    .B1(_05486_),
    .B2(_05487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05488_));
 sky130_fd_sc_hd__nand4_2 _14587_ (.A(_05472_),
    .B(_05474_),
    .C(_05486_),
    .D(_05487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05489_));
 sky130_fd_sc_hd__a21o_2 _14588_ (.A1(_05486_),
    .A2(_05487_),
    .B1(_05476_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05490_));
 sky130_fd_sc_hd__o211ai_2 _14589_ (.A1(_05471_),
    .A2(_05473_),
    .B1(_05486_),
    .C1(_05487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05491_));
 sky130_fd_sc_hd__nand2_2 _14590_ (.A(_05312_),
    .B(_05319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05492_));
 sky130_fd_sc_hd__a21oi_2 _14591_ (.A1(_05313_),
    .A2(_05314_),
    .B1(_05311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05493_));
 sky130_fd_sc_hd__nand3_2 _14592_ (.A(_05488_),
    .B(_05492_),
    .C(_05489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05494_));
 sky130_fd_sc_hd__nand3_2 _14593_ (.A(_05490_),
    .B(_05491_),
    .C(_05493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_2 _14594_ (.A(_05353_),
    .B(_05358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05496_));
 sky130_fd_sc_hd__nand4_2 _14595_ (.A(_05353_),
    .B(_05358_),
    .C(_05494_),
    .D(_05495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05497_));
 sky130_fd_sc_hd__a22o_2 _14596_ (.A1(_05353_),
    .A2(_05358_),
    .B1(_05494_),
    .B2(_05495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05498_));
 sky130_fd_sc_hd__a21o_2 _14597_ (.A1(_05494_),
    .A2(_05495_),
    .B1(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05499_));
 sky130_fd_sc_hd__nand2_2 _14598_ (.A(_05495_),
    .B(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05500_));
 sky130_fd_sc_hd__nand3_2 _14599_ (.A(_05494_),
    .B(_05495_),
    .C(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05501_));
 sky130_fd_sc_hd__nand3_2 _14600_ (.A(_05465_),
    .B(_05497_),
    .C(_05498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05502_));
 sky130_fd_sc_hd__nand4_2 _14601_ (.A(_05463_),
    .B(_05464_),
    .C(_05499_),
    .D(_05501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05503_));
 sky130_fd_sc_hd__nand4_2 _14602_ (.A(_05463_),
    .B(_05464_),
    .C(_05497_),
    .D(_05498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05504_));
 sky130_fd_sc_hd__nand3_2 _14603_ (.A(_05465_),
    .B(_05499_),
    .C(_05501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05505_));
 sky130_fd_sc_hd__nand3_2 _14604_ (.A(_05414_),
    .B(_05502_),
    .C(_05503_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05506_));
 sky130_fd_sc_hd__nand3_2 _14605_ (.A(_05413_),
    .B(_05504_),
    .C(_05505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_2 _14606_ (.A(_05506_),
    .B(_05507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05508_));
 sky130_fd_sc_hd__nand2_2 _14607_ (.A(\b_l[15] ),
    .B(\a_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05509_));
 sky130_fd_sc_hd__o2bb2ai_2 _14608_ (.A1_N(_05334_),
    .A2_N(_05337_),
    .B1(_05361_),
    .B2(_05368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05510_));
 sky130_fd_sc_hd__and4_2 _14609_ (.A(_05334_),
    .B(_05337_),
    .C(_05362_),
    .D(_05369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05511_));
 sky130_fd_sc_hd__o2111ai_2 _14610_ (.A1(_01888_),
    .A2(_05044_),
    .B1(_05337_),
    .C1(_05362_),
    .D1(_05369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05512_));
 sky130_fd_sc_hd__and3_2 _14611_ (.A(_05509_),
    .B(_05510_),
    .C(_05512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05513_));
 sky130_fd_sc_hd__o211ai_2 _14612_ (.A1(_09384_),
    .A2(_09395_),
    .B1(_05510_),
    .C1(_05512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05514_));
 sky130_fd_sc_hd__a21oi_2 _14613_ (.A1(_05510_),
    .A2(_05512_),
    .B1(_05509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05515_));
 sky130_fd_sc_hd__a21o_2 _14614_ (.A1(_05510_),
    .A2(_05512_),
    .B1(_05509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_2 _14615_ (.A(_05514_),
    .B(_05516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05517_));
 sky130_fd_sc_hd__nor2_2 _14616_ (.A(_05513_),
    .B(_05515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05518_));
 sky130_fd_sc_hd__nand4_2 _14617_ (.A(_05506_),
    .B(_05507_),
    .C(_05514_),
    .D(_05516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05519_));
 sky130_fd_sc_hd__o2bb2ai_2 _14618_ (.A1_N(_05506_),
    .A2_N(_05507_),
    .B1(_05513_),
    .B2(_05515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05520_));
 sky130_fd_sc_hd__o211ai_2 _14619_ (.A1(_05513_),
    .A2(_05515_),
    .B1(_05506_),
    .C1(_05507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_2 _14620_ (.A(_05508_),
    .B(_05518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05522_));
 sky130_fd_sc_hd__nand3_2 _14621_ (.A(_05412_),
    .B(_05521_),
    .C(_05522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05523_));
 sky130_fd_sc_hd__nand3_2 _14622_ (.A(_05411_),
    .B(_05519_),
    .C(_05520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05524_));
 sky130_fd_sc_hd__and3_2 _14623_ (.A(_05385_),
    .B(\a_h[1] ),
    .C(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05525_));
 sky130_fd_sc_hd__a31o_2 _14624_ (.A1(\b_l[15] ),
    .A2(\a_h[1] ),
    .A3(_05385_),
    .B1(_05384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05526_));
 sky130_fd_sc_hd__a21oi_2 _14625_ (.A1(_05523_),
    .A2(_05524_),
    .B1(_05526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05527_));
 sky130_fd_sc_hd__a21o_2 _14626_ (.A1(_05523_),
    .A2(_05524_),
    .B1(_05526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05528_));
 sky130_fd_sc_hd__o211a_2 _14627_ (.A1(_05384_),
    .A2(_05525_),
    .B1(_05524_),
    .C1(_05523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05529_));
 sky130_fd_sc_hd__o211ai_2 _14628_ (.A1(_05384_),
    .A2(_05525_),
    .B1(_05524_),
    .C1(_05523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05530_));
 sky130_fd_sc_hd__o22a_2 _14629_ (.A1(_05395_),
    .A2(_05404_),
    .B1(_05527_),
    .B2(_05529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05531_));
 sky130_fd_sc_hd__o22ai_2 _14630_ (.A1(_05395_),
    .A2(_05404_),
    .B1(_05527_),
    .B2(_05529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05532_));
 sky130_fd_sc_hd__nand3_2 _14631_ (.A(_05405_),
    .B(_05528_),
    .C(_05530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05533_));
 sky130_fd_sc_hd__o21ai_2 _14632_ (.A1(_05406_),
    .A2(_05263_),
    .B1(_05408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05534_));
 sky130_fd_sc_hd__a21oi_2 _14633_ (.A1(_05532_),
    .A2(_05533_),
    .B1(_05534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05535_));
 sky130_fd_sc_hd__and3_2 _14634_ (.A(_05534_),
    .B(_05533_),
    .C(_05532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05536_));
 sky130_fd_sc_hd__nor3_2 _14635_ (.A(rst),
    .B(_05535_),
    .C(_05536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00323_));
 sky130_fd_sc_hd__a32oi_2 _14636_ (.A1(_05412_),
    .A2(_05521_),
    .A3(_05522_),
    .B1(_05524_),
    .B2(_05526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_2 _14637_ (.A1(_05509_),
    .A2(_05511_),
    .B1(_05510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05538_));
 sky130_fd_sc_hd__a31o_2 _14638_ (.A1(_05414_),
    .A2(_05502_),
    .A3(_05503_),
    .B1(_05517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05539_));
 sky130_fd_sc_hd__a21boi_2 _14639_ (.A1(_05507_),
    .A2(_05517_),
    .B1_N(_05506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05540_));
 sky130_fd_sc_hd__nor2_2 _14640_ (.A(_09384_),
    .B(_09406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05541_));
 sky130_fd_sc_hd__a31o_2 _14641_ (.A1(_05488_),
    .A2(_05492_),
    .A3(_05489_),
    .B1(_05496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05542_));
 sky130_fd_sc_hd__o211a_2 _14642_ (.A1(_05468_),
    .A2(_05471_),
    .B1(_05495_),
    .C1(_05542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05543_));
 sky130_fd_sc_hd__o211ai_2 _14643_ (.A1(_05468_),
    .A2(_05471_),
    .B1(_05495_),
    .C1(_05542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05544_));
 sky130_fd_sc_hd__o2111ai_2 _14644_ (.A1(_05333_),
    .A2(_05467_),
    .B1(_05472_),
    .C1(_05494_),
    .D1(_05500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05545_));
 sky130_fd_sc_hd__a21o_2 _14645_ (.A1(_05544_),
    .A2(_05545_),
    .B1(_05541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05546_));
 sky130_fd_sc_hd__and3_2 _14646_ (.A(_05544_),
    .B(_05545_),
    .C(_05541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05547_));
 sky130_fd_sc_hd__nand4_2 _14647_ (.A(_05544_),
    .B(_05545_),
    .C(\b_l[15] ),
    .D(\a_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05548_));
 sky130_fd_sc_hd__nand2_2 _14648_ (.A(_05546_),
    .B(_05548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05549_));
 sky130_fd_sc_hd__nand3_2 _14649_ (.A(_05464_),
    .B(_05497_),
    .C(_05498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_2 _14650_ (.A(_05463_),
    .B(_05550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_2 _14651_ (.A(\b_l[5] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05552_));
 sky130_fd_sc_hd__a22oi_2 _14652_ (.A1(\b_l[4] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05553_));
 sky130_fd_sc_hd__and4_2 _14653_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05554_));
 sky130_fd_sc_hd__nand4_2 _14654_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_2 _14655_ (.A1(_05553_),
    .A2(_05554_),
    .B1(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05556_));
 sky130_fd_sc_hd__a41o_2 _14656_ (.A1(\b_l[3] ),
    .A2(\b_l[4] ),
    .A3(\a_h[14] ),
    .A4(\a_h[15] ),
    .B1(_05552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05557_));
 sky130_fd_sc_hd__a211oi_2 _14657_ (.A1(\b_l[5] ),
    .A2(\a_h[13] ),
    .B1(_05553_),
    .C1(_05554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05558_));
 sky130_fd_sc_hd__o211a_2 _14658_ (.A1(_05553_),
    .A2(_05554_),
    .B1(\b_l[5] ),
    .C1(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05559_));
 sky130_fd_sc_hd__o21ai_2 _14659_ (.A1(_05553_),
    .A2(_05557_),
    .B1(_05556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05560_));
 sky130_fd_sc_hd__o2bb2ai_2 _14660_ (.A1_N(_05286_),
    .A2_N(_05452_),
    .B1(_05558_),
    .B2(_05559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05561_));
 sky130_fd_sc_hd__inv_2 _14661_ (.A(_05561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05562_));
 sky130_fd_sc_hd__o211ai_2 _14662_ (.A1(_04988_),
    .A2(_05285_),
    .B1(_05452_),
    .C1(_05560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_2 _14663_ (.A(_05561_),
    .B(_05563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05564_));
 sky130_fd_sc_hd__a21bo_2 _14664_ (.A1(_05418_),
    .A2(_05422_),
    .B1_N(_05421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05565_));
 sky130_fd_sc_hd__a21boi_2 _14665_ (.A1(_05418_),
    .A2(_05422_),
    .B1_N(_05421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05566_));
 sky130_fd_sc_hd__o22ai_2 _14666_ (.A1(_05271_),
    .A2(_05446_),
    .B1(_05441_),
    .B2(_05444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05567_));
 sky130_fd_sc_hd__o22a_2 _14667_ (.A1(_05271_),
    .A2(_05446_),
    .B1(_05441_),
    .B2(_05444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_2 _14668_ (.A(\b_l[8] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2_2 _14669_ (.A(\b_l[6] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_2 _14670_ (.A(\b_l[7] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05571_));
 sky130_fd_sc_hd__a22oi_2 _14671_ (.A1(\b_l[7] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_2 _14672_ (.A(_05570_),
    .B(_05571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05573_));
 sky130_fd_sc_hd__and4_2 _14673_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05574_));
 sky130_fd_sc_hd__nand4_2 _14674_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05575_));
 sky130_fd_sc_hd__o22ai_2 _14675_ (.A1(_09264_),
    .A2(_09482_),
    .B1(_05572_),
    .B2(_05574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05576_));
 sky130_fd_sc_hd__nand4_2 _14676_ (.A(_05573_),
    .B(_05575_),
    .C(\b_l[8] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05577_));
 sky130_fd_sc_hd__o211ai_2 _14677_ (.A1(_09264_),
    .A2(_09482_),
    .B1(_05573_),
    .C1(_05575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05578_));
 sky130_fd_sc_hd__a21o_2 _14678_ (.A1(_05573_),
    .A2(_05575_),
    .B1(_05569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05579_));
 sky130_fd_sc_hd__a21oi_2 _14679_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05580_));
 sky130_fd_sc_hd__nand3_2 _14680_ (.A(_05568_),
    .B(_05578_),
    .C(_05579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05581_));
 sky130_fd_sc_hd__a211o_2 _14681_ (.A1(_05576_),
    .A2(_05577_),
    .B1(_05566_),
    .C1(_05567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05582_));
 sky130_fd_sc_hd__nand3_2 _14682_ (.A(_05576_),
    .B(_05577_),
    .C(_05567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05583_));
 sky130_fd_sc_hd__a31oi_2 _14683_ (.A1(_05576_),
    .A2(_05577_),
    .A3(_05567_),
    .B1(_05566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05584_));
 sky130_fd_sc_hd__a32oi_2 _14684_ (.A1(_05568_),
    .A2(_05578_),
    .A3(_05579_),
    .B1(_05583_),
    .B2(_05565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05585_));
 sky130_fd_sc_hd__o21ai_2 _14685_ (.A1(_05580_),
    .A2(_05584_),
    .B1(_05582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05586_));
 sky130_fd_sc_hd__a21o_2 _14686_ (.A1(_05581_),
    .A2(_05583_),
    .B1(_05566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05587_));
 sky130_fd_sc_hd__nand3_2 _14687_ (.A(_05566_),
    .B(_05581_),
    .C(_05583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05588_));
 sky130_fd_sc_hd__o211ai_2 _14688_ (.A1(_05565_),
    .A2(_05583_),
    .B1(_05586_),
    .C1(_05564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05589_));
 sky130_fd_sc_hd__nand4_2 _14689_ (.A(_05561_),
    .B(_05563_),
    .C(_05587_),
    .D(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05590_));
 sky130_fd_sc_hd__nand3_2 _14690_ (.A(_05564_),
    .B(_05587_),
    .C(_05588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05591_));
 sky130_fd_sc_hd__o2111ai_2 _14691_ (.A1(_05583_),
    .A2(_05565_),
    .B1(_05563_),
    .C1(_05561_),
    .D1(_05586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_2 _14692_ (.A(_05589_),
    .B(_05590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05593_));
 sky130_fd_sc_hd__nand3_2 _14693_ (.A(_05433_),
    .B(_05434_),
    .C(_05456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_2 _14694_ (.A(_05458_),
    .B(_05594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05595_));
 sky130_fd_sc_hd__nand3_2 _14695_ (.A(_05595_),
    .B(_05592_),
    .C(_05591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05596_));
 sky130_fd_sc_hd__nor2_2 _14696_ (.A(_05595_),
    .B(_05593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05597_));
 sky130_fd_sc_hd__nand4_2 _14697_ (.A(_05458_),
    .B(_05589_),
    .C(_05590_),
    .D(_05594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05598_));
 sky130_fd_sc_hd__a21bo_2 _14698_ (.A1(_05475_),
    .A2(_05486_),
    .B1_N(_05487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05599_));
 sky130_fd_sc_hd__a32oi_2 _14699_ (.A1(_05417_),
    .A2(_05423_),
    .A3(_05425_),
    .B1(_05428_),
    .B2(_05432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05600_));
 sky130_fd_sc_hd__o2bb2ai_2 _14700_ (.A1_N(_05432_),
    .A2_N(_05428_),
    .B1(_05424_),
    .B2(_05429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05601_));
 sky130_fd_sc_hd__nand2_2 _14701_ (.A(\b_l[12] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05602_));
 sky130_fd_sc_hd__nand2_2 _14702_ (.A(_05466_),
    .B(_05602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05603_));
 sky130_fd_sc_hd__nand2_2 _14703_ (.A(\b_l[13] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05604_));
 sky130_fd_sc_hd__nand4_2 _14704_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[5] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05605_));
 sky130_fd_sc_hd__o2111ai_2 _14705_ (.A1(_05467_),
    .A2(_05604_),
    .B1(\b_l[14] ),
    .C1(\a_h[4] ),
    .D1(_05603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05606_));
 sky130_fd_sc_hd__a22o_2 _14706_ (.A1(\b_l[14] ),
    .A2(\a_h[4] ),
    .B1(_05603_),
    .B2(_05605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05607_));
 sky130_fd_sc_hd__nand2_2 _14707_ (.A(_05606_),
    .B(_05607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05608_));
 sky130_fd_sc_hd__nand2_2 _14708_ (.A(_05478_),
    .B(_05481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_2 _14709_ (.A(_05480_),
    .B(_05609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05610_));
 sky130_fd_sc_hd__a21boi_2 _14710_ (.A1(_05478_),
    .A2(_05481_),
    .B1_N(_05480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05611_));
 sky130_fd_sc_hd__nand2_2 _14711_ (.A(\b_l[11] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05612_));
 sky130_fd_sc_hd__nand2_2 _14712_ (.A(\b_l[10] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05613_));
 sky130_fd_sc_hd__nand2_2 _14713_ (.A(\b_l[9] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05614_));
 sky130_fd_sc_hd__a22o_2 _14714_ (.A1(\b_l[10] ),
    .A2(\a_h[8] ),
    .B1(\a_h[9] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05615_));
 sky130_fd_sc_hd__nand2_2 _14715_ (.A(\b_l[10] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05616_));
 sky130_fd_sc_hd__nand4_2 _14716_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05617_));
 sky130_fd_sc_hd__o2bb2ai_2 _14717_ (.A1_N(_05613_),
    .A2_N(_05614_),
    .B1(_05616_),
    .B2(_05479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05618_));
 sky130_fd_sc_hd__o21ai_2 _14718_ (.A1(_09308_),
    .A2(_09449_),
    .B1(_05618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05619_));
 sky130_fd_sc_hd__o2111ai_2 _14719_ (.A1(_05479_),
    .A2(_05616_),
    .B1(\b_l[11] ),
    .C1(\a_h[7] ),
    .D1(_05615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05620_));
 sky130_fd_sc_hd__and3_2 _14720_ (.A(_05611_),
    .B(_05619_),
    .C(_05620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05621_));
 sky130_fd_sc_hd__nand3_2 _14721_ (.A(_05611_),
    .B(_05619_),
    .C(_05620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05622_));
 sky130_fd_sc_hd__o221ai_2 _14722_ (.A1(_09308_),
    .A2(_09449_),
    .B1(_05479_),
    .B2(_05616_),
    .C1(_05615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05623_));
 sky130_fd_sc_hd__nand3_2 _14723_ (.A(_05618_),
    .B(\a_h[7] ),
    .C(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05624_));
 sky130_fd_sc_hd__nand3_2 _14724_ (.A(_05624_),
    .B(_05610_),
    .C(_05623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05625_));
 sky130_fd_sc_hd__and3_2 _14725_ (.A(_05606_),
    .B(_05607_),
    .C(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05626_));
 sky130_fd_sc_hd__nand4_2 _14726_ (.A(_05606_),
    .B(_05607_),
    .C(_05622_),
    .D(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05627_));
 sky130_fd_sc_hd__a22o_2 _14727_ (.A1(_05606_),
    .A2(_05607_),
    .B1(_05622_),
    .B2(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05628_));
 sky130_fd_sc_hd__nand3_2 _14728_ (.A(_05628_),
    .B(_05600_),
    .C(_05627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_2 _14729_ (.A(_05608_),
    .B(_05625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05630_));
 sky130_fd_sc_hd__a21o_2 _14730_ (.A1(_05622_),
    .A2(_05625_),
    .B1(_05608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05631_));
 sky130_fd_sc_hd__o211ai_2 _14731_ (.A1(_05630_),
    .A2(_05621_),
    .B1(_05601_),
    .C1(_05631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05632_));
 sky130_fd_sc_hd__a31o_2 _14732_ (.A1(_05600_),
    .A2(_05627_),
    .A3(_05628_),
    .B1(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05633_));
 sky130_fd_sc_hd__nand2_2 _14733_ (.A(_05632_),
    .B(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05634_));
 sky130_fd_sc_hd__a21oi_2 _14734_ (.A1(_05629_),
    .A2(_05632_),
    .B1(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05635_));
 sky130_fd_sc_hd__a21o_2 _14735_ (.A1(_05629_),
    .A2(_05632_),
    .B1(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05636_));
 sky130_fd_sc_hd__and3_2 _14736_ (.A(_05629_),
    .B(_05632_),
    .C(_05599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05637_));
 sky130_fd_sc_hd__nand3_2 _14737_ (.A(_05632_),
    .B(_05599_),
    .C(_05629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05638_));
 sky130_fd_sc_hd__o2bb2ai_2 _14738_ (.A1_N(_05596_),
    .A2_N(_05598_),
    .B1(_05635_),
    .B2(_05637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05639_));
 sky130_fd_sc_hd__nand4_2 _14739_ (.A(_05596_),
    .B(_05598_),
    .C(_05636_),
    .D(_05638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_2 _14740_ (.A(_05639_),
    .B(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05641_));
 sky130_fd_sc_hd__and4_2 _14741_ (.A(_05463_),
    .B(_05550_),
    .C(_05639_),
    .D(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05642_));
 sky130_fd_sc_hd__nand4_2 _14742_ (.A(_05463_),
    .B(_05550_),
    .C(_05639_),
    .D(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05643_));
 sky130_fd_sc_hd__a22oi_2 _14743_ (.A1(_05463_),
    .A2(_05550_),
    .B1(_05639_),
    .B2(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05644_));
 sky130_fd_sc_hd__a22o_2 _14744_ (.A1(_05463_),
    .A2(_05550_),
    .B1(_05639_),
    .B2(_05640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05645_));
 sky130_fd_sc_hd__a21oi_2 _14745_ (.A1(_05641_),
    .A2(_05551_),
    .B1(_05549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05646_));
 sky130_fd_sc_hd__a21o_2 _14746_ (.A1(_05551_),
    .A2(_05641_),
    .B1(_05549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05647_));
 sky130_fd_sc_hd__a22o_2 _14747_ (.A1(_05546_),
    .A2(_05548_),
    .B1(_05643_),
    .B2(_05645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05648_));
 sky130_fd_sc_hd__o2111ai_2 _14748_ (.A1(_05647_),
    .A2(_05642_),
    .B1(_05539_),
    .C1(_05507_),
    .D1(_05648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05649_));
 sky130_fd_sc_hd__a22o_2 _14749_ (.A1(_05546_),
    .A2(_05548_),
    .B1(_05641_),
    .B2(_05551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05650_));
 sky130_fd_sc_hd__a21o_2 _14750_ (.A1(_05643_),
    .A2(_05645_),
    .B1(_05549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05651_));
 sky130_fd_sc_hd__o211ai_2 _14751_ (.A1(_05650_),
    .A2(_05642_),
    .B1(_05540_),
    .C1(_05651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05652_));
 sky130_fd_sc_hd__a21bo_2 _14752_ (.A1(_05649_),
    .A2(_05652_),
    .B1_N(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05653_));
 sky130_fd_sc_hd__o2111ai_2 _14753_ (.A1(_05511_),
    .A2(_05509_),
    .B1(_05510_),
    .C1(_05649_),
    .D1(_05652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_2 _14754_ (.A(_05652_),
    .B(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05655_));
 sky130_fd_sc_hd__nand3_2 _14755_ (.A(_05649_),
    .B(_05652_),
    .C(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05656_));
 sky130_fd_sc_hd__a21o_2 _14756_ (.A1(_05649_),
    .A2(_05652_),
    .B1(_05538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05657_));
 sky130_fd_sc_hd__nand3b_2 _14757_ (.A_N(_05537_),
    .B(_05656_),
    .C(_05657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05658_));
 sky130_fd_sc_hd__nand3_2 _14758_ (.A(_05653_),
    .B(_05654_),
    .C(_05537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_2 _14759_ (.A(_05658_),
    .B(_05659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05660_));
 sky130_fd_sc_hd__and4_2 _14760_ (.A(_05407_),
    .B(_05408_),
    .C(_05532_),
    .D(_05533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05661_));
 sky130_fd_sc_hd__nand4_2 _14761_ (.A(_05407_),
    .B(_05408_),
    .C(_05532_),
    .D(_05533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05662_));
 sky130_fd_sc_hd__nand3_2 _14762_ (.A(_05262_),
    .B(_05661_),
    .C(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05663_));
 sky130_fd_sc_hd__a21o_2 _14763_ (.A1(_05408_),
    .A2(_05533_),
    .B1(_05531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05664_));
 sky130_fd_sc_hd__o211ai_2 _14764_ (.A1(_05263_),
    .A2(_05662_),
    .B1(_05664_),
    .C1(_05660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05665_));
 sky130_fd_sc_hd__a21o_2 _14765_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05666_));
 sky130_fd_sc_hd__and3_2 _14766_ (.A(_09690_),
    .B(_05665_),
    .C(_05666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00324_));
 sky130_fd_sc_hd__a31o_2 _14767_ (.A1(\b_l[15] ),
    .A2(\a_h[3] ),
    .A3(_05545_),
    .B1(_05543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05667_));
 sky130_fd_sc_hd__nand3_2 _14768_ (.A(_05596_),
    .B(_05636_),
    .C(_05638_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05668_));
 sky130_fd_sc_hd__a31oi_2 _14769_ (.A1(_05596_),
    .A2(_05636_),
    .A3(_05638_),
    .B1(_05597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_2 _14770_ (.A(_05598_),
    .B(_05668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05670_));
 sky130_fd_sc_hd__o211ai_2 _14771_ (.A1(_05583_),
    .A2(_05565_),
    .B1(_05561_),
    .C1(_05586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05671_));
 sky130_fd_sc_hd__a31oi_2 _14772_ (.A1(_05563_),
    .A2(_05587_),
    .A3(_05588_),
    .B1(_05562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05672_));
 sky130_fd_sc_hd__and2_2 _14773_ (.A(\b_l[5] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05673_));
 sky130_fd_sc_hd__nand2_2 _14774_ (.A(\b_l[5] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05674_));
 sky130_fd_sc_hd__and4_2 _14775_ (.A(\b_l[4] ),
    .B(\b_l[5] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05675_));
 sky130_fd_sc_hd__a22oi_2 _14776_ (.A1(\b_l[5] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05676_));
 sky130_fd_sc_hd__nor2_2 _14777_ (.A(_05675_),
    .B(_05676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05677_));
 sky130_fd_sc_hd__a21o_2 _14778_ (.A1(_05552_),
    .A2(_05555_),
    .B1(_05553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05678_));
 sky130_fd_sc_hd__a21oi_2 _14779_ (.A1(_05552_),
    .A2(_05555_),
    .B1(_05553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_2 _14780_ (.A(\b_l[8] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05680_));
 sky130_fd_sc_hd__nand2_2 _14781_ (.A(\b_l[6] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_2 _14782_ (.A(\b_l[7] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_2 _14783_ (.A(_05681_),
    .B(_05682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05683_));
 sky130_fd_sc_hd__and4_2 _14784_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05684_));
 sky130_fd_sc_hd__nand4_2 _14785_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05685_));
 sky130_fd_sc_hd__a21bo_2 _14786_ (.A1(_05683_),
    .A2(_05685_),
    .B1_N(_05680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05686_));
 sky130_fd_sc_hd__nand4_2 _14787_ (.A(_05683_),
    .B(_05685_),
    .C(\b_l[8] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05687_));
 sky130_fd_sc_hd__o211ai_2 _14788_ (.A1(_09264_),
    .A2(_09493_),
    .B1(_05683_),
    .C1(_05685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05688_));
 sky130_fd_sc_hd__a21o_2 _14789_ (.A1(_05683_),
    .A2(_05685_),
    .B1(_05680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05689_));
 sky130_fd_sc_hd__nand2_2 _14790_ (.A(_05686_),
    .B(_05687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05690_));
 sky130_fd_sc_hd__and3_2 _14791_ (.A(_05689_),
    .B(_05678_),
    .C(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05691_));
 sky130_fd_sc_hd__nand3_2 _14792_ (.A(_05689_),
    .B(_05678_),
    .C(_05688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05692_));
 sky130_fd_sc_hd__nand3_2 _14793_ (.A(_05679_),
    .B(_05686_),
    .C(_05687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05693_));
 sky130_fd_sc_hd__o32a_2 _14794_ (.A1(_09493_),
    .A2(_09504_),
    .A3(_04260_),
    .B1(_09482_),
    .B2(_09264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05694_));
 sky130_fd_sc_hd__and3_2 _14795_ (.A(_05573_),
    .B(\a_h[10] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05695_));
 sky130_fd_sc_hd__a31o_2 _14796_ (.A1(\b_l[8] ),
    .A2(_05573_),
    .A3(\a_h[10] ),
    .B1(_05574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05696_));
 sky130_fd_sc_hd__o211ai_2 _14797_ (.A1(_05574_),
    .A2(_05695_),
    .B1(_05693_),
    .C1(_05692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05697_));
 sky130_fd_sc_hd__o2bb2ai_2 _14798_ (.A1_N(_05692_),
    .A2_N(_05693_),
    .B1(_05694_),
    .B2(_05572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05698_));
 sky130_fd_sc_hd__o2bb2ai_2 _14799_ (.A1_N(_05692_),
    .A2_N(_05693_),
    .B1(_05695_),
    .B2(_05574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05699_));
 sky130_fd_sc_hd__o2111ai_2 _14800_ (.A1(_05569_),
    .A2(_05572_),
    .B1(_05575_),
    .C1(_05692_),
    .D1(_05693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05700_));
 sky130_fd_sc_hd__and3_2 _14801_ (.A(_05698_),
    .B(_05677_),
    .C(_05697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05701_));
 sky130_fd_sc_hd__nand3_2 _14802_ (.A(_05698_),
    .B(_05677_),
    .C(_05697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05702_));
 sky130_fd_sc_hd__nand3b_2 _14803_ (.A_N(_05677_),
    .B(_05699_),
    .C(_05700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_2 _14804_ (.A(_05702_),
    .B(_05703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05704_));
 sky130_fd_sc_hd__nor2_2 _14805_ (.A(_05704_),
    .B(_05672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05705_));
 sky130_fd_sc_hd__nand4_2 _14806_ (.A(_05563_),
    .B(_05671_),
    .C(_05702_),
    .D(_05703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_2 _14807_ (.A(_05672_),
    .B(_05704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05707_));
 sky130_fd_sc_hd__nand2_2 _14808_ (.A(_05706_),
    .B(_05707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_2 _14809_ (.A(\b_l[12] ),
    .B(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05709_));
 sky130_fd_sc_hd__nand4_2 _14810_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[6] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_2 _14811_ (.A(_05604_),
    .B(_05709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05711_));
 sky130_fd_sc_hd__nand4_2 _14812_ (.A(_05711_),
    .B(\a_h[5] ),
    .C(\b_l[14] ),
    .D(_05710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05712_));
 sky130_fd_sc_hd__a22o_2 _14813_ (.A1(\b_l[14] ),
    .A2(\a_h[5] ),
    .B1(_05710_),
    .B2(_05711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05713_));
 sky130_fd_sc_hd__nand2_2 _14814_ (.A(_05712_),
    .B(_05713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_2 _14815_ (.A(\b_l[11] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05715_));
 sky130_fd_sc_hd__nand2_2 _14816_ (.A(\b_l[9] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05716_));
 sky130_fd_sc_hd__a22oi_2 _14817_ (.A1(\b_l[10] ),
    .A2(\a_h[9] ),
    .B1(\a_h[10] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_2 _14818_ (.A(_05616_),
    .B(_05716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05718_));
 sky130_fd_sc_hd__nand4_2 _14819_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05719_));
 sky130_fd_sc_hd__a21o_2 _14820_ (.A1(_05718_),
    .A2(_05719_),
    .B1(_05715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05720_));
 sky130_fd_sc_hd__o211ai_2 _14821_ (.A1(_09308_),
    .A2(_09460_),
    .B1(_05718_),
    .C1(_05719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05721_));
 sky130_fd_sc_hd__o2bb2ai_2 _14822_ (.A1_N(_05718_),
    .A2_N(_05719_),
    .B1(_09308_),
    .B2(_09460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05722_));
 sky130_fd_sc_hd__nand4_2 _14823_ (.A(_05718_),
    .B(_05719_),
    .C(\b_l[11] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05723_));
 sky130_fd_sc_hd__a22o_2 _14824_ (.A1(_05613_),
    .A2(_05614_),
    .B1(_05617_),
    .B2(_05612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05724_));
 sky130_fd_sc_hd__a22oi_2 _14825_ (.A1(_05613_),
    .A2(_05614_),
    .B1(_05617_),
    .B2(_05612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05725_));
 sky130_fd_sc_hd__nand3_2 _14826_ (.A(_05720_),
    .B(_05721_),
    .C(_05724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05726_));
 sky130_fd_sc_hd__nand3_2 _14827_ (.A(_05722_),
    .B(_05723_),
    .C(_05725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05727_));
 sky130_fd_sc_hd__a21oi_2 _14828_ (.A1(_05726_),
    .A2(_05727_),
    .B1(_05714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05728_));
 sky130_fd_sc_hd__a21o_2 _14829_ (.A1(_05726_),
    .A2(_05727_),
    .B1(_05714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05729_));
 sky130_fd_sc_hd__nand3_2 _14830_ (.A(_05714_),
    .B(_05726_),
    .C(_05727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05730_));
 sky130_fd_sc_hd__a22o_2 _14831_ (.A1(_05712_),
    .A2(_05713_),
    .B1(_05726_),
    .B2(_05727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05731_));
 sky130_fd_sc_hd__nand4_2 _14832_ (.A(_05712_),
    .B(_05713_),
    .C(_05726_),
    .D(_05727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05732_));
 sky130_fd_sc_hd__nand3_2 _14833_ (.A(_05731_),
    .B(_05732_),
    .C(_05585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_2 _14834_ (.A1(_05580_),
    .A2(_05584_),
    .B1(_05730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05734_));
 sky130_fd_sc_hd__o2111ai_2 _14835_ (.A1(_05565_),
    .A2(_05580_),
    .B1(_05583_),
    .C1(_05729_),
    .D1(_05730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05735_));
 sky130_fd_sc_hd__a31o_2 _14836_ (.A1(_05606_),
    .A2(_05607_),
    .A3(_05625_),
    .B1(_05621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05736_));
 sky130_fd_sc_hd__inv_2 _14837_ (.A(_05736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05737_));
 sky130_fd_sc_hd__o21ai_2 _14838_ (.A1(_05728_),
    .A2(_05734_),
    .B1(_05736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05738_));
 sky130_fd_sc_hd__o21ai_2 _14839_ (.A1(_05728_),
    .A2(_05734_),
    .B1(_05733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05739_));
 sky130_fd_sc_hd__o221a_2 _14840_ (.A1(_05621_),
    .A2(_05626_),
    .B1(_05728_),
    .B2(_05734_),
    .C1(_05733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05740_));
 sky130_fd_sc_hd__o221ai_2 _14841_ (.A1(_05621_),
    .A2(_05626_),
    .B1(_05728_),
    .B2(_05734_),
    .C1(_05733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05741_));
 sky130_fd_sc_hd__a21oi_2 _14842_ (.A1(_05733_),
    .A2(_05735_),
    .B1(_05736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05742_));
 sky130_fd_sc_hd__nand2_2 _14843_ (.A(_05739_),
    .B(_05737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05743_));
 sky130_fd_sc_hd__o21ai_2 _14844_ (.A1(_05740_),
    .A2(_05742_),
    .B1(_05708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05744_));
 sky130_fd_sc_hd__nand4_2 _14845_ (.A(_05706_),
    .B(_05707_),
    .C(_05741_),
    .D(_05743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05745_));
 sky130_fd_sc_hd__nand3_2 _14846_ (.A(_05708_),
    .B(_05741_),
    .C(_05743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05746_));
 sky130_fd_sc_hd__o211ai_2 _14847_ (.A1(_05740_),
    .A2(_05742_),
    .B1(_05706_),
    .C1(_05707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05747_));
 sky130_fd_sc_hd__a21oi_2 _14848_ (.A1(_05744_),
    .A2(_05745_),
    .B1(_05670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05748_));
 sky130_fd_sc_hd__nand3_2 _14849_ (.A(_05669_),
    .B(_05746_),
    .C(_05747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05749_));
 sky130_fd_sc_hd__a21oi_2 _14850_ (.A1(_05746_),
    .A2(_05747_),
    .B1(_05669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05750_));
 sky130_fd_sc_hd__nand3_2 _14851_ (.A(_05670_),
    .B(_05744_),
    .C(_05745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05751_));
 sky130_fd_sc_hd__nand2_2 _14852_ (.A(_05749_),
    .B(_05751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05752_));
 sky130_fd_sc_hd__o21ai_2 _14853_ (.A1(_05467_),
    .A2(_05604_),
    .B1(_05606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05753_));
 sky130_fd_sc_hd__nand3_2 _14854_ (.A(_05632_),
    .B(_05633_),
    .C(_05753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05754_));
 sky130_fd_sc_hd__o2111ai_2 _14855_ (.A1(_05467_),
    .A2(_05604_),
    .B1(_05606_),
    .C1(_05629_),
    .D1(_05634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05755_));
 sky130_fd_sc_hd__inv_2 _14856_ (.A(_05755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05756_));
 sky130_fd_sc_hd__nand2_2 _14857_ (.A(\b_l[15] ),
    .B(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05757_));
 sky130_fd_sc_hd__a32o_2 _14858_ (.A1(_05632_),
    .A2(_05633_),
    .A3(_05753_),
    .B1(\a_h[4] ),
    .B2(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05758_));
 sky130_fd_sc_hd__a21o_2 _14859_ (.A1(_05754_),
    .A2(_05755_),
    .B1(_05757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05759_));
 sky130_fd_sc_hd__nand4_2 _14860_ (.A(_05754_),
    .B(_05755_),
    .C(\b_l[15] ),
    .D(\a_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05760_));
 sky130_fd_sc_hd__a22o_2 _14861_ (.A1(\b_l[15] ),
    .A2(\a_h[4] ),
    .B1(_05754_),
    .B2(_05755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05761_));
 sky130_fd_sc_hd__o21a_2 _14862_ (.A1(_05756_),
    .A2(_05758_),
    .B1(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05762_));
 sky130_fd_sc_hd__o21ai_2 _14863_ (.A1(_05756_),
    .A2(_05758_),
    .B1(_05759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05763_));
 sky130_fd_sc_hd__nand4_2 _14864_ (.A(_05749_),
    .B(_05751_),
    .C(_05760_),
    .D(_05761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05764_));
 sky130_fd_sc_hd__nand2_2 _14865_ (.A(_05752_),
    .B(_05762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05765_));
 sky130_fd_sc_hd__o2111ai_2 _14866_ (.A1(_05756_),
    .A2(_05758_),
    .B1(_05759_),
    .C1(_05751_),
    .D1(_05749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_2 _14867_ (.A1(_05748_),
    .A2(_05750_),
    .B1(_05763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05767_));
 sky130_fd_sc_hd__o21a_2 _14868_ (.A1(_05549_),
    .A2(_05644_),
    .B1(_05643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05768_));
 sky130_fd_sc_hd__nand3_2 _14869_ (.A(_05768_),
    .B(_05767_),
    .C(_05766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05769_));
 sky130_fd_sc_hd__o211ai_2 _14870_ (.A1(_05642_),
    .A2(_05646_),
    .B1(_05764_),
    .C1(_05765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05770_));
 sky130_fd_sc_hd__a21oi_2 _14871_ (.A1(_05769_),
    .A2(_05770_),
    .B1(_05667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05771_));
 sky130_fd_sc_hd__o211a_2 _14872_ (.A1(_05543_),
    .A2(_05547_),
    .B1(_05769_),
    .C1(_05770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05772_));
 sky130_fd_sc_hd__o211ai_2 _14873_ (.A1(_05543_),
    .A2(_05547_),
    .B1(_05769_),
    .C1(_05770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05773_));
 sky130_fd_sc_hd__nand2_2 _14874_ (.A(_05649_),
    .B(_05655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05774_));
 sky130_fd_sc_hd__nand3b_2 _14875_ (.A_N(_05771_),
    .B(_05774_),
    .C(_05773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05775_));
 sky130_fd_sc_hd__o211a_2 _14876_ (.A1(_05771_),
    .A2(_05772_),
    .B1(_05649_),
    .C1(_05655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05776_));
 sky130_fd_sc_hd__o211ai_2 _14877_ (.A1(_05771_),
    .A2(_05772_),
    .B1(_05649_),
    .C1(_05655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_2 _14878_ (.A(_05775_),
    .B(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05778_));
 sky130_fd_sc_hd__a21oi_2 _14879_ (.A1(_05658_),
    .A2(_05666_),
    .B1(_05778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05779_));
 sky130_fd_sc_hd__a31o_2 _14880_ (.A1(_05658_),
    .A2(_05666_),
    .A3(_05778_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05780_));
 sky130_fd_sc_hd__nor2_2 _14881_ (.A(_05779_),
    .B(_05780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00325_));
 sky130_fd_sc_hd__a21boi_2 _14882_ (.A1(_05667_),
    .A2(_05769_),
    .B1_N(_05770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05781_));
 sky130_fd_sc_hd__a32oi_2 _14883_ (.A1(_05670_),
    .A2(_05744_),
    .A3(_05745_),
    .B1(_05760_),
    .B2(_05761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05782_));
 sky130_fd_sc_hd__a31o_2 _14884_ (.A1(_05749_),
    .A2(_05760_),
    .A3(_05761_),
    .B1(_05750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05783_));
 sky130_fd_sc_hd__o2111a_2 _14885_ (.A1(_05604_),
    .A2(_05709_),
    .B1(_05712_),
    .C1(_05733_),
    .D1(_05738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05784_));
 sky130_fd_sc_hd__o2111ai_2 _14886_ (.A1(_05604_),
    .A2(_05709_),
    .B1(_05712_),
    .C1(_05733_),
    .D1(_05738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05785_));
 sky130_fd_sc_hd__a22oi_2 _14887_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05733_),
    .B2(_05738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05786_));
 sky130_fd_sc_hd__a22o_2 _14888_ (.A1(_05710_),
    .A2(_05712_),
    .B1(_05733_),
    .B2(_05738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05787_));
 sky130_fd_sc_hd__nor2_2 _14889_ (.A(_09384_),
    .B(_09428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_2 _14890_ (.A1(_05784_),
    .A2(_05786_),
    .B1(_05788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05789_));
 sky130_fd_sc_hd__o211ai_2 _14891_ (.A1(_09384_),
    .A2(_09428_),
    .B1(_05785_),
    .C1(_05787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_2 _14892_ (.A(_05789_),
    .B(_05790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05791_));
 sky130_fd_sc_hd__a31oi_2 _14893_ (.A1(_05707_),
    .A2(_05741_),
    .A3(_05743_),
    .B1(_05705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05792_));
 sky130_fd_sc_hd__a31o_2 _14894_ (.A1(_05707_),
    .A2(_05741_),
    .A3(_05743_),
    .B1(_05705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05793_));
 sky130_fd_sc_hd__nand2_2 _14895_ (.A(\b_l[6] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05794_));
 sky130_fd_sc_hd__nand2_2 _14896_ (.A(\b_l[7] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_2 _14897_ (.A(_05794_),
    .B(_05795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05796_));
 sky130_fd_sc_hd__nand2_2 _14898_ (.A(\b_l[7] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05797_));
 sky130_fd_sc_hd__and4_2 _14899_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[13] ),
    .D(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05798_));
 sky130_fd_sc_hd__nand4_2 _14900_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[13] ),
    .D(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05799_));
 sky130_fd_sc_hd__and2_2 _14901_ (.A(\b_l[8] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05800_));
 sky130_fd_sc_hd__a21oi_2 _14902_ (.A1(_05796_),
    .A2(_05799_),
    .B1(_05800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05801_));
 sky130_fd_sc_hd__o2bb2ai_2 _14903_ (.A1_N(_05796_),
    .A2_N(_05799_),
    .B1(_09264_),
    .B2(_09504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05802_));
 sky130_fd_sc_hd__o211a_2 _14904_ (.A1(_05681_),
    .A2(_05797_),
    .B1(_05800_),
    .C1(_05796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05803_));
 sky130_fd_sc_hd__o2111ai_2 _14905_ (.A1(_05681_),
    .A2(_05797_),
    .B1(\b_l[8] ),
    .C1(\a_h[12] ),
    .D1(_05796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05804_));
 sky130_fd_sc_hd__nor2_2 _14906_ (.A(_05801_),
    .B(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05805_));
 sky130_fd_sc_hd__nand3_2 _14907_ (.A(_05802_),
    .B(_05804_),
    .C(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05806_));
 sky130_fd_sc_hd__a21oi_2 _14908_ (.A1(_05802_),
    .A2(_05804_),
    .B1(_05675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05807_));
 sky130_fd_sc_hd__o22ai_2 _14909_ (.A1(_05446_),
    .A2(_05674_),
    .B1(_05801_),
    .B2(_05803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05808_));
 sky130_fd_sc_hd__a31o_2 _14910_ (.A1(\b_l[8] ),
    .A2(_05683_),
    .A3(\a_h[11] ),
    .B1(_05684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05809_));
 sky130_fd_sc_hd__a31oi_2 _14911_ (.A1(_05683_),
    .A2(\a_h[11] ),
    .A3(\b_l[8] ),
    .B1(_05684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05810_));
 sky130_fd_sc_hd__a21oi_2 _14912_ (.A1(_05806_),
    .A2(_05808_),
    .B1(_05809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05811_));
 sky130_fd_sc_hd__a21o_2 _14913_ (.A1(_05806_),
    .A2(_05808_),
    .B1(_05809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05812_));
 sky130_fd_sc_hd__nand3_2 _14914_ (.A(_05806_),
    .B(_05808_),
    .C(_05809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05813_));
 sky130_fd_sc_hd__and3_2 _14915_ (.A(_05806_),
    .B(_05808_),
    .C(_05810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05814_));
 sky130_fd_sc_hd__o21ai_2 _14916_ (.A1(_05810_),
    .A2(_05805_),
    .B1(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05815_));
 sky130_fd_sc_hd__a31o_2 _14917_ (.A1(_05806_),
    .A2(_05808_),
    .A3(_05809_),
    .B1(_05674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05816_));
 sky130_fd_sc_hd__nand4_2 _14918_ (.A(_05812_),
    .B(_05813_),
    .C(\b_l[5] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05817_));
 sky130_fd_sc_hd__o22ai_2 _14919_ (.A1(_05815_),
    .A2(_05814_),
    .B1(_05811_),
    .B2(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_2 _14920_ (.A(_05702_),
    .B(_05818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05819_));
 sky130_fd_sc_hd__o211ai_2 _14921_ (.A1(_05814_),
    .A2(_05815_),
    .B1(_05817_),
    .C1(_05701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_2 _14922_ (.A(\b_l[10] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2_2 _14923_ (.A(\b_l[9] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05822_));
 sky130_fd_sc_hd__a22oi_2 _14924_ (.A1(\b_l[10] ),
    .A2(\a_h[10] ),
    .B1(\a_h[11] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2_2 _14925_ (.A(_05821_),
    .B(_05822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05824_));
 sky130_fd_sc_hd__nand4_2 _14926_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_2 _14927_ (.A(\b_l[11] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05826_));
 sky130_fd_sc_hd__a21bo_2 _14928_ (.A1(_05824_),
    .A2(_05825_),
    .B1_N(_05826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05827_));
 sky130_fd_sc_hd__a41o_2 _14929_ (.A1(\b_l[9] ),
    .A2(\b_l[10] ),
    .A3(\a_h[10] ),
    .A4(\a_h[11] ),
    .B1(_05826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05828_));
 sky130_fd_sc_hd__a21o_2 _14930_ (.A1(_05824_),
    .A2(_05825_),
    .B1(_05826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05829_));
 sky130_fd_sc_hd__o211ai_2 _14931_ (.A1(_09308_),
    .A2(_09471_),
    .B1(_05824_),
    .C1(_05825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05830_));
 sky130_fd_sc_hd__o21a_2 _14932_ (.A1(_05616_),
    .A2(_05716_),
    .B1(_05715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05831_));
 sky130_fd_sc_hd__a21oi_2 _14933_ (.A1(_05715_),
    .A2(_05719_),
    .B1(_05717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05832_));
 sky130_fd_sc_hd__o211ai_2 _14934_ (.A1(_05717_),
    .A2(_05831_),
    .B1(_05830_),
    .C1(_05829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05833_));
 sky130_fd_sc_hd__o211ai_2 _14935_ (.A1(_05823_),
    .A2(_05828_),
    .B1(_05832_),
    .C1(_05827_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05834_));
 sky130_fd_sc_hd__nand2_2 _14936_ (.A(\b_l[14] ),
    .B(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05835_));
 sky130_fd_sc_hd__a22oi_2 _14937_ (.A1(\b_l[13] ),
    .A2(\a_h[7] ),
    .B1(\a_h[8] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05836_));
 sky130_fd_sc_hd__a22o_2 _14938_ (.A1(\b_l[13] ),
    .A2(\a_h[7] ),
    .B1(\a_h[8] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05837_));
 sky130_fd_sc_hd__and4_2 _14939_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05838_));
 sky130_fd_sc_hd__nand4_2 _14940_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[7] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05839_));
 sky130_fd_sc_hd__and4_2 _14941_ (.A(_05837_),
    .B(_05839_),
    .C(\b_l[14] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05840_));
 sky130_fd_sc_hd__o22a_2 _14942_ (.A1(_09362_),
    .A2(_09439_),
    .B1(_05836_),
    .B2(_05838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05841_));
 sky130_fd_sc_hd__o211a_2 _14943_ (.A1(_05836_),
    .A2(_05838_),
    .B1(\b_l[14] ),
    .C1(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05842_));
 sky130_fd_sc_hd__o311a_2 _14944_ (.A1(_09449_),
    .A2(_09460_),
    .A3(_05044_),
    .B1(_05835_),
    .C1(_05837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05843_));
 sky130_fd_sc_hd__nor2_2 _14945_ (.A(_05840_),
    .B(_05841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05844_));
 sky130_fd_sc_hd__o2bb2ai_2 _14946_ (.A1_N(_05833_),
    .A2_N(_05834_),
    .B1(_05840_),
    .B2(_05841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05845_));
 sky130_fd_sc_hd__nand3_2 _14947_ (.A(_05844_),
    .B(_05834_),
    .C(_05833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05846_));
 sky130_fd_sc_hd__a31oi_2 _14948_ (.A1(_05679_),
    .A2(_05686_),
    .A3(_05687_),
    .B1(_05696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05847_));
 sky130_fd_sc_hd__nand2_2 _14949_ (.A(_05692_),
    .B(_05696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05848_));
 sky130_fd_sc_hd__o21ai_2 _14950_ (.A1(_05678_),
    .A2(_05690_),
    .B1(_05848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05849_));
 sky130_fd_sc_hd__nand3_2 _14951_ (.A(_05845_),
    .B(_05846_),
    .C(_05849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05850_));
 sky130_fd_sc_hd__o211ai_2 _14952_ (.A1(_05840_),
    .A2(_05841_),
    .B1(_05833_),
    .C1(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05851_));
 sky130_fd_sc_hd__o2bb2ai_2 _14953_ (.A1_N(_05833_),
    .A2_N(_05834_),
    .B1(_05842_),
    .B2(_05843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05852_));
 sky130_fd_sc_hd__o211ai_2 _14954_ (.A1(_05691_),
    .A2(_05847_),
    .B1(_05851_),
    .C1(_05852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05853_));
 sky130_fd_sc_hd__nand2_2 _14955_ (.A(_05850_),
    .B(_05853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05854_));
 sky130_fd_sc_hd__a21bo_2 _14956_ (.A1(_05714_),
    .A2(_05727_),
    .B1_N(_05726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05855_));
 sky130_fd_sc_hd__a21boi_2 _14957_ (.A1(_05714_),
    .A2(_05727_),
    .B1_N(_05726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_2 _14958_ (.A(_05854_),
    .B(_05856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05857_));
 sky130_fd_sc_hd__nand3_2 _14959_ (.A(_05850_),
    .B(_05853_),
    .C(_05855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05858_));
 sky130_fd_sc_hd__nand3_2 _14960_ (.A(_05850_),
    .B(_05853_),
    .C(_05856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05859_));
 sky130_fd_sc_hd__a21o_2 _14961_ (.A1(_05850_),
    .A2(_05853_),
    .B1(_05856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05860_));
 sky130_fd_sc_hd__a22o_2 _14962_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_05859_),
    .B2(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05861_));
 sky130_fd_sc_hd__nand4_2 _14963_ (.A(_05819_),
    .B(_05820_),
    .C(_05859_),
    .D(_05860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05862_));
 sky130_fd_sc_hd__nand4_2 _14964_ (.A(_05819_),
    .B(_05820_),
    .C(_05857_),
    .D(_05858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05863_));
 sky130_fd_sc_hd__a22o_2 _14965_ (.A1(_05819_),
    .A2(_05820_),
    .B1(_05857_),
    .B2(_05858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05864_));
 sky130_fd_sc_hd__nand2_2 _14966_ (.A(_05861_),
    .B(_05862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05865_));
 sky130_fd_sc_hd__and3_2 _14967_ (.A(_05793_),
    .B(_05861_),
    .C(_05862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05866_));
 sky130_fd_sc_hd__nand3_2 _14968_ (.A(_05793_),
    .B(_05861_),
    .C(_05862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05867_));
 sky130_fd_sc_hd__nand3_2 _14969_ (.A(_05864_),
    .B(_05792_),
    .C(_05863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05868_));
 sky130_fd_sc_hd__nand4_2 _14970_ (.A(_05789_),
    .B(_05790_),
    .C(_05867_),
    .D(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05869_));
 sky130_fd_sc_hd__a22o_2 _14971_ (.A1(_05789_),
    .A2(_05790_),
    .B1(_05867_),
    .B2(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05870_));
 sky130_fd_sc_hd__nand2_2 _14972_ (.A(_05791_),
    .B(_05868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05871_));
 sky130_fd_sc_hd__a21o_2 _14973_ (.A1(_05867_),
    .A2(_05868_),
    .B1(_05791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05872_));
 sky130_fd_sc_hd__o211ai_2 _14974_ (.A1(_05866_),
    .A2(_05871_),
    .B1(_05872_),
    .C1(_05783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05873_));
 sky130_fd_sc_hd__o211ai_2 _14975_ (.A1(_05748_),
    .A2(_05782_),
    .B1(_05869_),
    .C1(_05870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05874_));
 sky130_fd_sc_hd__o31a_2 _14976_ (.A1(_09384_),
    .A2(_09417_),
    .A3(_05756_),
    .B1(_05754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05875_));
 sky130_fd_sc_hd__inv_2 _14977_ (.A(_05875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05876_));
 sky130_fd_sc_hd__a21o_2 _14978_ (.A1(_05873_),
    .A2(_05874_),
    .B1(_05875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05877_));
 sky130_fd_sc_hd__o2111ai_2 _14979_ (.A1(_05757_),
    .A2(_05756_),
    .B1(_05754_),
    .C1(_05874_),
    .D1(_05873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05878_));
 sky130_fd_sc_hd__nand4_2 _14980_ (.A(_05755_),
    .B(_05758_),
    .C(_05873_),
    .D(_05874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05879_));
 sky130_fd_sc_hd__a22o_2 _14981_ (.A1(_05755_),
    .A2(_05758_),
    .B1(_05873_),
    .B2(_05874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05880_));
 sky130_fd_sc_hd__nand4_2 _14982_ (.A(_05770_),
    .B(_05773_),
    .C(_05877_),
    .D(_05878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05881_));
 sky130_fd_sc_hd__a21oi_2 _14983_ (.A1(_05877_),
    .A2(_05878_),
    .B1(_05781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05882_));
 sky130_fd_sc_hd__nand3b_2 _14984_ (.A_N(_05781_),
    .B(_05879_),
    .C(_05880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05883_));
 sky130_fd_sc_hd__nand2_2 _14985_ (.A(_05881_),
    .B(_05883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05884_));
 sky130_fd_sc_hd__a21o_2 _14986_ (.A1(_05658_),
    .A2(_05775_),
    .B1(_05776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05885_));
 sky130_fd_sc_hd__nand4_2 _14987_ (.A(_05658_),
    .B(_05659_),
    .C(_05775_),
    .D(_05777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05886_));
 sky130_fd_sc_hd__nor2_2 _14988_ (.A(_05662_),
    .B(_05886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05887_));
 sky130_fd_sc_hd__nand3_2 _14989_ (.A(_05262_),
    .B(_05887_),
    .C(_05260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05888_));
 sky130_fd_sc_hd__o21a_2 _14990_ (.A1(_05886_),
    .A2(_05664_),
    .B1(_05885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05889_));
 sky130_fd_sc_hd__o21ai_2 _14991_ (.A1(_05663_),
    .A2(_05886_),
    .B1(_05889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05890_));
 sky130_fd_sc_hd__and2_2 _14992_ (.A(_05889_),
    .B(_05884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05891_));
 sky130_fd_sc_hd__and3_2 _14993_ (.A(_05890_),
    .B(_05883_),
    .C(_05881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05892_));
 sky130_fd_sc_hd__a211oi_2 _14994_ (.A1(_05891_),
    .A2(_05888_),
    .B1(rst),
    .C1(_05892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00326_));
 sky130_fd_sc_hd__a21boi_2 _14995_ (.A1(_05874_),
    .A2(_05876_),
    .B1_N(_05873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_2 _14996_ (.A1(_05792_),
    .A2(_05865_),
    .B1(_05871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_2 _14997_ (.A(_05853_),
    .B(_05856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05895_));
 sky130_fd_sc_hd__o2111ai_2 _14998_ (.A1(_05835_),
    .A2(_05836_),
    .B1(_05839_),
    .C1(_05850_),
    .D1(_05895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05896_));
 sky130_fd_sc_hd__inv_2 _14999_ (.A(_05896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_2 _15000_ (.A(_05850_),
    .B(_05855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05898_));
 sky130_fd_sc_hd__o211ai_2 _15001_ (.A1(_05838_),
    .A2(_05840_),
    .B1(_05853_),
    .C1(_05898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05899_));
 sky130_fd_sc_hd__a22o_2 _15002_ (.A1(\b_l[15] ),
    .A2(\a_h[6] ),
    .B1(_05896_),
    .B2(_05899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05900_));
 sky130_fd_sc_hd__nand4_2 _15003_ (.A(_05896_),
    .B(_05899_),
    .C(\b_l[15] ),
    .D(\a_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05901_));
 sky130_fd_sc_hd__nand2_2 _15004_ (.A(_05900_),
    .B(_05901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05902_));
 sky130_fd_sc_hd__nand3_2 _15005_ (.A(_05820_),
    .B(_05857_),
    .C(_05858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_2 _15006_ (.A(_05819_),
    .B(_05903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05904_));
 sky130_fd_sc_hd__a31o_2 _15007_ (.A1(\b_l[8] ),
    .A2(_05796_),
    .A3(\a_h[12] ),
    .B1(_05798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05905_));
 sky130_fd_sc_hd__nand2_2 _15008_ (.A(\b_l[6] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05906_));
 sky130_fd_sc_hd__nand4_2 _15009_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05907_));
 sky130_fd_sc_hd__nand2_2 _15010_ (.A(_05797_),
    .B(_05906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05908_));
 sky130_fd_sc_hd__a22o_2 _15011_ (.A1(\b_l[8] ),
    .A2(\a_h[13] ),
    .B1(_05907_),
    .B2(_05908_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05909_));
 sky130_fd_sc_hd__nand4_2 _15012_ (.A(_05908_),
    .B(\a_h[13] ),
    .C(\b_l[8] ),
    .D(_05907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05910_));
 sky130_fd_sc_hd__a21oi_2 _15013_ (.A1(_05909_),
    .A2(_05910_),
    .B1(_05905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05911_));
 sky130_fd_sc_hd__and3_2 _15014_ (.A(_05905_),
    .B(_05909_),
    .C(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05912_));
 sky130_fd_sc_hd__o211ai_2 _15015_ (.A1(_05798_),
    .A2(_05803_),
    .B1(_05909_),
    .C1(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05913_));
 sky130_fd_sc_hd__nor2_2 _15016_ (.A(_05911_),
    .B(_05912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05914_));
 sky130_fd_sc_hd__o22a_2 _15017_ (.A1(_05911_),
    .A2(_05912_),
    .B1(_05811_),
    .B2(_05816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05915_));
 sky130_fd_sc_hd__a31o_2 _15018_ (.A1(_05812_),
    .A2(_05813_),
    .A3(_05673_),
    .B1(_05914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05916_));
 sky130_fd_sc_hd__and4_2 _15019_ (.A(_05812_),
    .B(_05914_),
    .C(_05813_),
    .D(_05673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05917_));
 sky130_fd_sc_hd__nand4_2 _15020_ (.A(_05812_),
    .B(_05914_),
    .C(_05813_),
    .D(_05673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05918_));
 sky130_fd_sc_hd__a21bo_2 _15021_ (.A1(_05844_),
    .A2(_05833_),
    .B1_N(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05919_));
 sky130_fd_sc_hd__a21boi_2 _15022_ (.A1(_05844_),
    .A2(_05833_),
    .B1_N(_05834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05920_));
 sky130_fd_sc_hd__a21boi_2 _15023_ (.A1(_05808_),
    .A2(_05809_),
    .B1_N(_05806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05921_));
 sky130_fd_sc_hd__o21ai_2 _15024_ (.A1(_05810_),
    .A2(_05807_),
    .B1(_05806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_2 _15025_ (.A(_05825_),
    .B(_05826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05923_));
 sky130_fd_sc_hd__o21ai_2 _15026_ (.A1(_05826_),
    .A2(_05823_),
    .B1(_05825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05924_));
 sky130_fd_sc_hd__nand2_2 _15027_ (.A(\b_l[11] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05925_));
 sky130_fd_sc_hd__nand2_2 _15028_ (.A(\b_l[9] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_2 _15029_ (.A(\b_l[10] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05927_));
 sky130_fd_sc_hd__nand4_2 _15030_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05928_));
 sky130_fd_sc_hd__a22oi_2 _15031_ (.A1(\b_l[10] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_2 _15032_ (.A(_05926_),
    .B(_05927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05930_));
 sky130_fd_sc_hd__o2bb2ai_2 _15033_ (.A1_N(_05928_),
    .A2_N(_05930_),
    .B1(_09308_),
    .B2(_09482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05931_));
 sky130_fd_sc_hd__nand4_2 _15034_ (.A(_05930_),
    .B(\a_h[10] ),
    .C(\b_l[11] ),
    .D(_05928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05932_));
 sky130_fd_sc_hd__a21oi_2 _15035_ (.A1(_05928_),
    .A2(_05930_),
    .B1(_05925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05933_));
 sky130_fd_sc_hd__nand2_2 _15036_ (.A(_05925_),
    .B(_05928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05934_));
 sky130_fd_sc_hd__o2bb2ai_2 _15037_ (.A1_N(_05824_),
    .A2_N(_05923_),
    .B1(_05929_),
    .B2(_05934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05935_));
 sky130_fd_sc_hd__a21oi_2 _15038_ (.A1(_05931_),
    .A2(_05932_),
    .B1(_05924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05936_));
 sky130_fd_sc_hd__nand3_2 _15039_ (.A(_05931_),
    .B(_05932_),
    .C(_05924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_2 _15040_ (.A1(_05933_),
    .A2(_05935_),
    .B1(_05937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05938_));
 sky130_fd_sc_hd__nand2_2 _15041_ (.A(\b_l[13] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05939_));
 sky130_fd_sc_hd__nand2_2 _15042_ (.A(\b_l[13] ),
    .B(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_2 _15043_ (.A(\b_l[12] ),
    .B(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05941_));
 sky130_fd_sc_hd__and4_2 _15044_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05942_));
 sky130_fd_sc_hd__nand4_2 _15045_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[8] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_2 _15046_ (.A(_05940_),
    .B(_05941_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05944_));
 sky130_fd_sc_hd__a22oi_2 _15047_ (.A1(\b_l[14] ),
    .A2(\a_h[7] ),
    .B1(_05943_),
    .B2(_05944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05945_));
 sky130_fd_sc_hd__a22o_2 _15048_ (.A1(\b_l[14] ),
    .A2(\a_h[7] ),
    .B1(_05943_),
    .B2(_05944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05946_));
 sky130_fd_sc_hd__and4_2 _15049_ (.A(_05944_),
    .B(\a_h[7] ),
    .C(\b_l[14] ),
    .D(_05943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05947_));
 sky130_fd_sc_hd__nand4_2 _15050_ (.A(_05944_),
    .B(\a_h[7] ),
    .C(\b_l[14] ),
    .D(_05943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05948_));
 sky130_fd_sc_hd__nor2_2 _15051_ (.A(_05945_),
    .B(_05947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05949_));
 sky130_fd_sc_hd__nand2_2 _15052_ (.A(_05946_),
    .B(_05948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05950_));
 sky130_fd_sc_hd__o21ai_2 _15053_ (.A1(_05945_),
    .A2(_05947_),
    .B1(_05938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05951_));
 sky130_fd_sc_hd__o211ai_2 _15054_ (.A1(_05933_),
    .A2(_05935_),
    .B1(_05937_),
    .C1(_05949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05952_));
 sky130_fd_sc_hd__o21ai_2 _15055_ (.A1(_05945_),
    .A2(_05947_),
    .B1(_05937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05953_));
 sky130_fd_sc_hd__nand2_2 _15056_ (.A(_05938_),
    .B(_05949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05954_));
 sky130_fd_sc_hd__nand3_2 _15057_ (.A(_05922_),
    .B(_05951_),
    .C(_05952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05955_));
 sky130_fd_sc_hd__inv_2 _15058_ (.A(_05955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05956_));
 sky130_fd_sc_hd__o211ai_2 _15059_ (.A1(_05936_),
    .A2(_05953_),
    .B1(_05954_),
    .C1(_05921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05957_));
 sky130_fd_sc_hd__a21o_2 _15060_ (.A1(_05955_),
    .A2(_05957_),
    .B1(_05919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05958_));
 sky130_fd_sc_hd__nand2_2 _15061_ (.A(_05957_),
    .B(_05919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05959_));
 sky130_fd_sc_hd__nand3_2 _15062_ (.A(_05920_),
    .B(_05955_),
    .C(_05957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05960_));
 sky130_fd_sc_hd__a21o_2 _15063_ (.A1(_05955_),
    .A2(_05957_),
    .B1(_05920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05961_));
 sky130_fd_sc_hd__nand3_2 _15064_ (.A(_05918_),
    .B(_05960_),
    .C(_05961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05962_));
 sky130_fd_sc_hd__nand4_2 _15065_ (.A(_05916_),
    .B(_05918_),
    .C(_05960_),
    .D(_05961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05963_));
 sky130_fd_sc_hd__o221ai_2 _15066_ (.A1(_05956_),
    .A2(_05959_),
    .B1(_05915_),
    .B2(_05917_),
    .C1(_05958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05964_));
 sky130_fd_sc_hd__o2111ai_2 _15067_ (.A1(_05959_),
    .A2(_05956_),
    .B1(_05918_),
    .C1(_05916_),
    .D1(_05958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05965_));
 sky130_fd_sc_hd__o211ai_2 _15068_ (.A1(_05915_),
    .A2(_05917_),
    .B1(_05960_),
    .C1(_05961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05966_));
 sky130_fd_sc_hd__a21oi_2 _15069_ (.A1(_05963_),
    .A2(_05964_),
    .B1(_05904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05967_));
 sky130_fd_sc_hd__nand4_2 _15070_ (.A(_05819_),
    .B(_05903_),
    .C(_05965_),
    .D(_05966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05968_));
 sky130_fd_sc_hd__a22oi_2 _15071_ (.A1(_05819_),
    .A2(_05903_),
    .B1(_05965_),
    .B2(_05966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05969_));
 sky130_fd_sc_hd__a22o_2 _15072_ (.A1(_05819_),
    .A2(_05903_),
    .B1(_05965_),
    .B2(_05966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05970_));
 sky130_fd_sc_hd__a21oi_2 _15073_ (.A1(_05968_),
    .A2(_05970_),
    .B1(_05902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05971_));
 sky130_fd_sc_hd__nand3_2 _15074_ (.A(_05970_),
    .B(_05902_),
    .C(_05968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05972_));
 sky130_fd_sc_hd__nand4_2 _15075_ (.A(_05900_),
    .B(_05901_),
    .C(_05968_),
    .D(_05970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05973_));
 sky130_fd_sc_hd__o21ai_2 _15076_ (.A1(_05967_),
    .A2(_05969_),
    .B1(_05902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05974_));
 sky130_fd_sc_hd__nand3_2 _15077_ (.A(_05894_),
    .B(_05973_),
    .C(_05974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05975_));
 sky130_fd_sc_hd__o211ai_2 _15078_ (.A1(_05792_),
    .A2(_05865_),
    .B1(_05871_),
    .C1(_05972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05976_));
 sky130_fd_sc_hd__o21ai_2 _15079_ (.A1(_05971_),
    .A2(_05976_),
    .B1(_05975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05977_));
 sky130_fd_sc_hd__a31o_2 _15080_ (.A1(_05785_),
    .A2(\a_h[5] ),
    .A3(\b_l[15] ),
    .B1(_05786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05978_));
 sky130_fd_sc_hd__o31a_2 _15081_ (.A1(_09384_),
    .A2(_09428_),
    .A3(_05784_),
    .B1(_05787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05979_));
 sky130_fd_sc_hd__o211ai_2 _15082_ (.A1(_05971_),
    .A2(_05976_),
    .B1(_05979_),
    .C1(_05975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05980_));
 sky130_fd_sc_hd__nand2_2 _15083_ (.A(_05977_),
    .B(_05978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05981_));
 sky130_fd_sc_hd__nand3_2 _15084_ (.A(_05893_),
    .B(_05980_),
    .C(_05981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05982_));
 sky130_fd_sc_hd__a21oi_2 _15085_ (.A1(_05980_),
    .A2(_05981_),
    .B1(_05893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05983_));
 sky130_fd_sc_hd__a21o_2 _15086_ (.A1(_05980_),
    .A2(_05981_),
    .B1(_05893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05984_));
 sky130_fd_sc_hd__nand2_2 _15087_ (.A(_05982_),
    .B(_05984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05985_));
 sky130_fd_sc_hd__a21oi_2 _15088_ (.A1(_05890_),
    .A2(_05881_),
    .B1(_05882_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05986_));
 sky130_fd_sc_hd__a21oi_2 _15089_ (.A1(_05986_),
    .A2(_05985_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05987_));
 sky130_fd_sc_hd__o21a_2 _15090_ (.A1(_05985_),
    .A2(_05986_),
    .B1(_05987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00327_));
 sky130_fd_sc_hd__a21o_2 _15091_ (.A1(_05902_),
    .A2(_05968_),
    .B1(_05969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05988_));
 sky130_fd_sc_hd__a21oi_2 _15092_ (.A1(_05902_),
    .A2(_05968_),
    .B1(_05969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05989_));
 sky130_fd_sc_hd__nand2_2 _15093_ (.A(_05920_),
    .B(_05955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05990_));
 sky130_fd_sc_hd__o211a_2 _15094_ (.A1(_05942_),
    .A2(_05947_),
    .B1(_05957_),
    .C1(_05990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05991_));
 sky130_fd_sc_hd__o211ai_2 _15095_ (.A1(_05942_),
    .A2(_05947_),
    .B1(_05957_),
    .C1(_05990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05992_));
 sky130_fd_sc_hd__o2111ai_2 _15096_ (.A1(_05940_),
    .A2(_05941_),
    .B1(_05948_),
    .C1(_05955_),
    .D1(_05959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05993_));
 sky130_fd_sc_hd__o2bb2ai_2 _15097_ (.A1_N(_05992_),
    .A2_N(_05993_),
    .B1(_09384_),
    .B2(_09449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05994_));
 sky130_fd_sc_hd__nand4_2 _15098_ (.A(_05992_),
    .B(_05993_),
    .C(\b_l[15] ),
    .D(\a_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05995_));
 sky130_fd_sc_hd__and2_2 _15099_ (.A(_05994_),
    .B(_05995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05996_));
 sky130_fd_sc_hd__nand2_2 _15100_ (.A(_05994_),
    .B(_05995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_05997_));
 sky130_fd_sc_hd__a31o_2 _15101_ (.A1(_05918_),
    .A2(_05960_),
    .A3(_05961_),
    .B1(_05915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05998_));
 sky130_fd_sc_hd__and4_2 _15102_ (.A(\b_l[7] ),
    .B(\b_l[8] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_05999_));
 sky130_fd_sc_hd__nand4_2 _15103_ (.A(\b_l[7] ),
    .B(\b_l[8] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06000_));
 sky130_fd_sc_hd__a22oi_2 _15104_ (.A1(\b_l[8] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06001_));
 sky130_fd_sc_hd__o221a_2 _15105_ (.A1(_05797_),
    .A2(_05906_),
    .B1(_05999_),
    .B2(_06001_),
    .C1(_05910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06002_));
 sky130_fd_sc_hd__a211oi_2 _15106_ (.A1(_05907_),
    .A2(_05910_),
    .B1(_05999_),
    .C1(_06001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06003_));
 sky130_fd_sc_hd__or2_2 _15107_ (.A(_06002_),
    .B(_06003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06004_));
 sky130_fd_sc_hd__o21a_2 _15108_ (.A1(_05950_),
    .A2(_05936_),
    .B1(_05937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06005_));
 sky130_fd_sc_hd__inv_2 _15109_ (.A(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_2 _15110_ (.A(\b_l[12] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06007_));
 sky130_fd_sc_hd__nand2_2 _15111_ (.A(_05939_),
    .B(_06007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_2 _15112_ (.A(\b_l[13] ),
    .B(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06009_));
 sky130_fd_sc_hd__and3_2 _15113_ (.A(\a_h[9] ),
    .B(\a_h[10] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06010_));
 sky130_fd_sc_hd__nand4_2 _15114_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[9] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06011_));
 sky130_fd_sc_hd__and4_2 _15115_ (.A(_06008_),
    .B(_06011_),
    .C(\b_l[14] ),
    .D(\a_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06012_));
 sky130_fd_sc_hd__or4b_2 _15116_ (.A(_09362_),
    .B(_06010_),
    .C(_09460_),
    .D_N(_06008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06013_));
 sky130_fd_sc_hd__a22oi_2 _15117_ (.A1(\b_l[14] ),
    .A2(\a_h[8] ),
    .B1(_06008_),
    .B2(_06011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06014_));
 sky130_fd_sc_hd__nor2_2 _15118_ (.A(_06012_),
    .B(_06014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06015_));
 sky130_fd_sc_hd__o21ai_2 _15119_ (.A1(_05925_),
    .A2(_05929_),
    .B1(_05928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06016_));
 sky130_fd_sc_hd__o21a_2 _15120_ (.A1(_05925_),
    .A2(_05929_),
    .B1(_05928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06017_));
 sky130_fd_sc_hd__nand2_2 _15121_ (.A(\b_l[11] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_2 _15122_ (.A(\b_l[9] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_2 _15123_ (.A(\b_l[10] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06020_));
 sky130_fd_sc_hd__nand4_2 _15124_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06021_));
 sky130_fd_sc_hd__a22oi_2 _15125_ (.A1(\b_l[10] ),
    .A2(\a_h[12] ),
    .B1(\a_h[13] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_2 _15126_ (.A(_06019_),
    .B(_06020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06023_));
 sky130_fd_sc_hd__o2bb2ai_2 _15127_ (.A1_N(_06021_),
    .A2_N(_06023_),
    .B1(_09308_),
    .B2(_09493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06024_));
 sky130_fd_sc_hd__nand4_2 _15128_ (.A(_06023_),
    .B(\a_h[11] ),
    .C(\b_l[11] ),
    .D(_06021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06025_));
 sky130_fd_sc_hd__a21oi_2 _15129_ (.A1(_06021_),
    .A2(_06023_),
    .B1(_06018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06026_));
 sky130_fd_sc_hd__a21o_2 _15130_ (.A1(_06021_),
    .A2(_06023_),
    .B1(_06018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06027_));
 sky130_fd_sc_hd__o21a_2 _15131_ (.A1(_06019_),
    .A2(_06020_),
    .B1(_06018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06028_));
 sky130_fd_sc_hd__o21ai_2 _15132_ (.A1(_06019_),
    .A2(_06020_),
    .B1(_06018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06029_));
 sky130_fd_sc_hd__o2bb2ai_2 _15133_ (.A1_N(_05930_),
    .A2_N(_05934_),
    .B1(_06022_),
    .B2(_06029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06030_));
 sky130_fd_sc_hd__o211ai_2 _15134_ (.A1(_06029_),
    .A2(_06022_),
    .B1(_06017_),
    .C1(_06027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06031_));
 sky130_fd_sc_hd__and3_2 _15135_ (.A(_06024_),
    .B(_06025_),
    .C(_06016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06032_));
 sky130_fd_sc_hd__nand3_2 _15136_ (.A(_06024_),
    .B(_06025_),
    .C(_06016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06033_));
 sky130_fd_sc_hd__o21ai_2 _15137_ (.A1(_06026_),
    .A2(_06030_),
    .B1(_06033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06034_));
 sky130_fd_sc_hd__o211ai_2 _15138_ (.A1(_06012_),
    .A2(_06014_),
    .B1(_06031_),
    .C1(_06033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06035_));
 sky130_fd_sc_hd__nand2_2 _15139_ (.A(_06034_),
    .B(_06015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06036_));
 sky130_fd_sc_hd__nand3_2 _15140_ (.A(_05913_),
    .B(_06035_),
    .C(_06036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06037_));
 sky130_fd_sc_hd__o211ai_2 _15141_ (.A1(_06026_),
    .A2(_06030_),
    .B1(_06033_),
    .C1(_06015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_2 _15142_ (.A1(_06012_),
    .A2(_06014_),
    .B1(_06034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06039_));
 sky130_fd_sc_hd__nand3_2 _15143_ (.A(_06039_),
    .B(_05912_),
    .C(_06038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06040_));
 sky130_fd_sc_hd__nand2_2 _15144_ (.A(_06040_),
    .B(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06041_));
 sky130_fd_sc_hd__nand3_2 _15145_ (.A(_06037_),
    .B(_06040_),
    .C(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06042_));
 sky130_fd_sc_hd__a21o_2 _15146_ (.A1(_06037_),
    .A2(_06040_),
    .B1(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06043_));
 sky130_fd_sc_hd__nand3_2 _15147_ (.A(_06006_),
    .B(_06037_),
    .C(_06040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06044_));
 sky130_fd_sc_hd__a21o_2 _15148_ (.A1(_06037_),
    .A2(_06040_),
    .B1(_06006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06045_));
 sky130_fd_sc_hd__o211ai_2 _15149_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_06042_),
    .C1(_06043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06046_));
 sky130_fd_sc_hd__nand3b_2 _15150_ (.A_N(_06004_),
    .B(_06044_),
    .C(_06045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06047_));
 sky130_fd_sc_hd__nand2_2 _15151_ (.A(_06046_),
    .B(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06048_));
 sky130_fd_sc_hd__and4_2 _15152_ (.A(_05916_),
    .B(_05962_),
    .C(_06046_),
    .D(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06049_));
 sky130_fd_sc_hd__nand4_2 _15153_ (.A(_05916_),
    .B(_05962_),
    .C(_06046_),
    .D(_06047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_2 _15154_ (.A(_05998_),
    .B(_06048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06051_));
 sky130_fd_sc_hd__nand3_2 _15155_ (.A(_05997_),
    .B(_06050_),
    .C(_06051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06052_));
 sky130_fd_sc_hd__a21o_2 _15156_ (.A1(_06050_),
    .A2(_06051_),
    .B1(_05997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06053_));
 sky130_fd_sc_hd__a21oi_2 _15157_ (.A1(_05998_),
    .A2(_06048_),
    .B1(_05997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06054_));
 sky130_fd_sc_hd__a21o_2 _15158_ (.A1(_05998_),
    .A2(_06048_),
    .B1(_05997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06055_));
 sky130_fd_sc_hd__and3_2 _15159_ (.A(_05996_),
    .B(_06050_),
    .C(_06051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06056_));
 sky130_fd_sc_hd__a22o_2 _15160_ (.A1(_05994_),
    .A2(_05995_),
    .B1(_06050_),
    .B2(_06051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06057_));
 sky130_fd_sc_hd__nand3_2 _15161_ (.A(_06053_),
    .B(_05988_),
    .C(_06052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_2 _15162_ (.A(_05989_),
    .B(_06057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06059_));
 sky130_fd_sc_hd__o211ai_2 _15163_ (.A1(_06055_),
    .A2(_06049_),
    .B1(_05989_),
    .C1(_06057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_2 _15164_ (.A(_06058_),
    .B(_06060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06061_));
 sky130_fd_sc_hd__o21a_2 _15165_ (.A1(_09384_),
    .A2(_09439_),
    .B1(_05899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06062_));
 sky130_fd_sc_hd__nor2_2 _15166_ (.A(_05897_),
    .B(_06062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_2 _15167_ (.A(_06061_),
    .B(_06063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06064_));
 sky130_fd_sc_hd__o211ai_2 _15168_ (.A1(_05897_),
    .A2(_06062_),
    .B1(_06060_),
    .C1(_06058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06065_));
 sky130_fd_sc_hd__o2bb2ai_2 _15169_ (.A1_N(_06058_),
    .A2_N(_06060_),
    .B1(_06062_),
    .B2(_05897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06066_));
 sky130_fd_sc_hd__nand3_2 _15170_ (.A(_06058_),
    .B(_06060_),
    .C(_06063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06067_));
 sky130_fd_sc_hd__a2bb2oi_2 _15171_ (.A1_N(_05971_),
    .A2_N(_05976_),
    .B1(_05979_),
    .B2(_05975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06068_));
 sky130_fd_sc_hd__o2bb2ai_2 _15172_ (.A1_N(_05975_),
    .A2_N(_05979_),
    .B1(_05976_),
    .B2(_05971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06069_));
 sky130_fd_sc_hd__nand3_2 _15173_ (.A(_06064_),
    .B(_06065_),
    .C(_06069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06070_));
 sky130_fd_sc_hd__and3_2 _15174_ (.A(_06066_),
    .B(_06067_),
    .C(_06068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06071_));
 sky130_fd_sc_hd__nand3_2 _15175_ (.A(_06066_),
    .B(_06067_),
    .C(_06068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_2 _15176_ (.A(_06070_),
    .B(_06072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06073_));
 sky130_fd_sc_hd__a21o_2 _15177_ (.A1(_05882_),
    .A2(_05982_),
    .B1(_05983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06074_));
 sky130_fd_sc_hd__nor2_2 _15178_ (.A(_05884_),
    .B(_05985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06075_));
 sky130_fd_sc_hd__a21boi_2 _15179_ (.A1(_05888_),
    .A2(_05889_),
    .B1_N(_06075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06076_));
 sky130_fd_sc_hd__a221oi_2 _15180_ (.A1(_06070_),
    .A2(_06072_),
    .B1(_06075_),
    .B2(_05890_),
    .C1(_06074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06077_));
 sky130_fd_sc_hd__o21bai_2 _15181_ (.A1(_06074_),
    .A2(_06076_),
    .B1_N(_06073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06078_));
 sky130_fd_sc_hd__nor3b_2 _15182_ (.A(rst),
    .B(_06077_),
    .C_N(_06078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00328_));
 sky130_fd_sc_hd__o2bb2ai_2 _15183_ (.A1_N(_06063_),
    .A2_N(_06058_),
    .B1(_06056_),
    .B2(_06059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06079_));
 sky130_fd_sc_hd__a31o_2 _15184_ (.A1(\b_l[15] ),
    .A2(_05993_),
    .A3(\a_h[7] ),
    .B1(_05991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06080_));
 sky130_fd_sc_hd__inv_2 _15185_ (.A(_06080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06081_));
 sky130_fd_sc_hd__a21oi_2 _15186_ (.A1(_05996_),
    .A2(_06051_),
    .B1(_06049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06082_));
 sky130_fd_sc_hd__nor2_2 _15187_ (.A(_09384_),
    .B(_09460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06083_));
 sky130_fd_sc_hd__a31o_2 _15188_ (.A1(_05913_),
    .A2(_06035_),
    .A3(_06036_),
    .B1(_06005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06084_));
 sky130_fd_sc_hd__o211ai_2 _15189_ (.A1(_06010_),
    .A2(_06012_),
    .B1(_06037_),
    .C1(_06041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06085_));
 sky130_fd_sc_hd__o2111ai_2 _15190_ (.A1(_02278_),
    .A2(_05044_),
    .B1(_06013_),
    .C1(_06040_),
    .D1(_06084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06086_));
 sky130_fd_sc_hd__a21oi_2 _15191_ (.A1(_06085_),
    .A2(_06086_),
    .B1(_06083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06087_));
 sky130_fd_sc_hd__and3_2 _15192_ (.A(_06086_),
    .B(_06083_),
    .C(_06085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06088_));
 sky130_fd_sc_hd__nor2_2 _15193_ (.A(_06087_),
    .B(_06088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06089_));
 sky130_fd_sc_hd__and3_2 _15194_ (.A(_05797_),
    .B(\a_h[15] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06090_));
 sky130_fd_sc_hd__nand2_2 _15195_ (.A(\b_l[9] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_2 _15196_ (.A(\b_l[10] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06092_));
 sky130_fd_sc_hd__a22oi_2 _15197_ (.A1(\b_l[10] ),
    .A2(\a_h[13] ),
    .B1(\a_h[14] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06093_));
 sky130_fd_sc_hd__nand2_2 _15198_ (.A(_06091_),
    .B(_06092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_2 _15199_ (.A(\b_l[10] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06095_));
 sky130_fd_sc_hd__nand4_2 _15200_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[13] ),
    .D(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06096_));
 sky130_fd_sc_hd__o2bb2ai_2 _15201_ (.A1_N(_06091_),
    .A2_N(_06092_),
    .B1(_06095_),
    .B2(_06019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06097_));
 sky130_fd_sc_hd__and2_2 _15202_ (.A(\b_l[11] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06098_));
 sky130_fd_sc_hd__nand2_2 _15203_ (.A(\b_l[11] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06099_));
 sky130_fd_sc_hd__nand3_2 _15204_ (.A(_06094_),
    .B(_06096_),
    .C(_06098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06100_));
 sky130_fd_sc_hd__a21oi_2 _15205_ (.A1(_06094_),
    .A2(_06096_),
    .B1(_06098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06101_));
 sky130_fd_sc_hd__o21ai_2 _15206_ (.A1(_09308_),
    .A2(_09504_),
    .B1(_06097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06102_));
 sky130_fd_sc_hd__a2bb2oi_2 _15207_ (.A1_N(_06022_),
    .A2_N(_06028_),
    .B1(_06100_),
    .B2(_06102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06103_));
 sky130_fd_sc_hd__a22o_2 _15208_ (.A1(_06023_),
    .A2(_06029_),
    .B1(_06100_),
    .B2(_06102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06104_));
 sky130_fd_sc_hd__nand3_2 _15209_ (.A(_06023_),
    .B(_06029_),
    .C(_06100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06105_));
 sky130_fd_sc_hd__nor2_2 _15210_ (.A(_06101_),
    .B(_06105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_2 _15211_ (.A(\b_l[12] ),
    .B(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06107_));
 sky130_fd_sc_hd__and3_2 _15212_ (.A(\a_h[10] ),
    .B(\a_h[11] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06108_));
 sky130_fd_sc_hd__nand4_2 _15213_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[10] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_2 _15214_ (.A(_06009_),
    .B(_06107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06110_));
 sky130_fd_sc_hd__a22oi_2 _15215_ (.A1(\b_l[14] ),
    .A2(\a_h[9] ),
    .B1(_06109_),
    .B2(_06110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06111_));
 sky130_fd_sc_hd__and4_2 _15216_ (.A(_06110_),
    .B(\a_h[9] ),
    .C(\b_l[14] ),
    .D(_06109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06112_));
 sky130_fd_sc_hd__nor2_2 _15217_ (.A(_06111_),
    .B(_06112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06113_));
 sky130_fd_sc_hd__o211ai_2 _15218_ (.A1(_06101_),
    .A2(_06105_),
    .B1(_06113_),
    .C1(_06104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06114_));
 sky130_fd_sc_hd__o21bai_2 _15219_ (.A1(_06103_),
    .A2(_06106_),
    .B1_N(_06113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06115_));
 sky130_fd_sc_hd__o221ai_2 _15220_ (.A1(_06101_),
    .A2(_06105_),
    .B1(_06111_),
    .B2(_06112_),
    .C1(_06104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06116_));
 sky130_fd_sc_hd__o21ai_2 _15221_ (.A1(_06103_),
    .A2(_06106_),
    .B1(_06113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06117_));
 sky130_fd_sc_hd__nand3b_2 _15222_ (.A_N(_06003_),
    .B(_06116_),
    .C(_06117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06118_));
 sky130_fd_sc_hd__nand3_2 _15223_ (.A(_06114_),
    .B(_06115_),
    .C(_06003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06119_));
 sky130_fd_sc_hd__o21ai_2 _15224_ (.A1(_06015_),
    .A2(_06032_),
    .B1(_06031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06120_));
 sky130_fd_sc_hd__o22a_2 _15225_ (.A1(_06030_),
    .A2(_06026_),
    .B1(_06015_),
    .B2(_06032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06121_));
 sky130_fd_sc_hd__a21o_2 _15226_ (.A1(_06118_),
    .A2(_06119_),
    .B1(_06121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06122_));
 sky130_fd_sc_hd__nand3_2 _15227_ (.A(_06118_),
    .B(_06119_),
    .C(_06121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06123_));
 sky130_fd_sc_hd__a21o_2 _15228_ (.A1(_06118_),
    .A2(_06119_),
    .B1(_06120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06124_));
 sky130_fd_sc_hd__nand3_2 _15229_ (.A(_06118_),
    .B(_06119_),
    .C(_06120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3b_2 _15230_ (.A_N(_06090_),
    .B(_06124_),
    .C(_06125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06126_));
 sky130_fd_sc_hd__nand3_2 _15231_ (.A(_06122_),
    .B(_06123_),
    .C(_06090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06127_));
 sky130_fd_sc_hd__nand2_2 _15232_ (.A(_06126_),
    .B(_06127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_2 _15233_ (.A(_06047_),
    .B(_06128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06129_));
 sky130_fd_sc_hd__nand3b_2 _15234_ (.A_N(_06047_),
    .B(_06126_),
    .C(_06127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2_2 _15235_ (.A(_06047_),
    .B(_06128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_2 _15236_ (.A(_06130_),
    .B(_06131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06132_));
 sky130_fd_sc_hd__nand2_2 _15237_ (.A(_06132_),
    .B(_06089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06133_));
 sky130_fd_sc_hd__o221ai_2 _15238_ (.A1(_06087_),
    .A2(_06088_),
    .B1(_06128_),
    .B2(_06047_),
    .C1(_06131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_2 _15239_ (.A(_06089_),
    .B(_06131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06135_));
 sky130_fd_sc_hd__a2bb2o_2 _15240_ (.A1_N(_06087_),
    .A2_N(_06088_),
    .B1(_06130_),
    .B2(_06131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06136_));
 sky130_fd_sc_hd__o221ai_2 _15241_ (.A1(_06049_),
    .A2(_06054_),
    .B1(_06129_),
    .B2(_06135_),
    .C1(_06136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06137_));
 sky130_fd_sc_hd__nand3_2 _15242_ (.A(_06082_),
    .B(_06133_),
    .C(_06134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06138_));
 sky130_fd_sc_hd__a21boi_2 _15243_ (.A1(_06080_),
    .A2(_06138_),
    .B1_N(_06137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06139_));
 sky130_fd_sc_hd__a21o_2 _15244_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06140_));
 sky130_fd_sc_hd__nand3_2 _15245_ (.A(_06137_),
    .B(_06138_),
    .C(_06080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06141_));
 sky130_fd_sc_hd__a21o_2 _15246_ (.A1(_06137_),
    .A2(_06138_),
    .B1(_06081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06142_));
 sky130_fd_sc_hd__nand3_2 _15247_ (.A(_06081_),
    .B(_06137_),
    .C(_06138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06143_));
 sky130_fd_sc_hd__nand3b_2 _15248_ (.A_N(_06079_),
    .B(_06142_),
    .C(_06143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06144_));
 sky130_fd_sc_hd__nand3_2 _15249_ (.A(_06140_),
    .B(_06141_),
    .C(_06079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_2 _15250_ (.A(_06144_),
    .B(_06145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06146_));
 sky130_fd_sc_hd__a21oi_2 _15251_ (.A1(_06072_),
    .A2(_06078_),
    .B1(_06146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06147_));
 sky130_fd_sc_hd__a31o_2 _15252_ (.A1(_06072_),
    .A2(_06078_),
    .A3(_06146_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06148_));
 sky130_fd_sc_hd__nor2_2 _15253_ (.A(_06147_),
    .B(_06148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00329_));
 sky130_fd_sc_hd__a22oi_2 _15254_ (.A1(\b_l[13] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06149_));
 sky130_fd_sc_hd__a22o_2 _15255_ (.A1(\b_l[13] ),
    .A2(\a_h[11] ),
    .B1(\a_h[12] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06150_));
 sky130_fd_sc_hd__and4_2 _15256_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06151_));
 sky130_fd_sc_hd__nand4_2 _15257_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[11] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06152_));
 sky130_fd_sc_hd__o22a_2 _15258_ (.A1(_09362_),
    .A2(_09482_),
    .B1(_06149_),
    .B2(_06151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06153_));
 sky130_fd_sc_hd__a22o_2 _15259_ (.A1(\b_l[14] ),
    .A2(\a_h[10] ),
    .B1(_06150_),
    .B2(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06154_));
 sky130_fd_sc_hd__and4_2 _15260_ (.A(_06150_),
    .B(_06152_),
    .C(\b_l[14] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06155_));
 sky130_fd_sc_hd__nand4_2 _15261_ (.A(_06150_),
    .B(_06152_),
    .C(\b_l[14] ),
    .D(\a_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06156_));
 sky130_fd_sc_hd__nor2_2 _15262_ (.A(_06153_),
    .B(_06155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_2 _15263_ (.A(_06154_),
    .B(_06156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06158_));
 sky130_fd_sc_hd__o21ai_2 _15264_ (.A1(_06099_),
    .A2(_06093_),
    .B1(_06096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06159_));
 sky130_fd_sc_hd__and2_2 _15265_ (.A(\b_l[11] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06160_));
 sky130_fd_sc_hd__nand2_2 _15266_ (.A(\b_l[11] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_2 _15267_ (.A(\b_l[10] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06162_));
 sky130_fd_sc_hd__nand4_2 _15268_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06163_));
 sky130_fd_sc_hd__nand2_2 _15269_ (.A(\b_l[9] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06164_));
 sky130_fd_sc_hd__a22oi_2 _15270_ (.A1(\b_l[10] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06165_));
 sky130_fd_sc_hd__nand2_2 _15271_ (.A(_06095_),
    .B(_06164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06166_));
 sky130_fd_sc_hd__o211a_2 _15272_ (.A1(_06091_),
    .A2(_06162_),
    .B1(_06160_),
    .C1(_06166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06167_));
 sky130_fd_sc_hd__o2111ai_2 _15273_ (.A1(_06091_),
    .A2(_06162_),
    .B1(\b_l[11] ),
    .C1(\a_h[13] ),
    .D1(_06166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06168_));
 sky130_fd_sc_hd__a21oi_2 _15274_ (.A1(_06163_),
    .A2(_06166_),
    .B1(_06160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06169_));
 sky130_fd_sc_hd__o2bb2ai_2 _15275_ (.A1_N(_06163_),
    .A2_N(_06166_),
    .B1(_09308_),
    .B2(_09515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06170_));
 sky130_fd_sc_hd__nand2_2 _15276_ (.A(_06159_),
    .B(_06170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06171_));
 sky130_fd_sc_hd__and3_2 _15277_ (.A(_06159_),
    .B(_06168_),
    .C(_06170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06172_));
 sky130_fd_sc_hd__nand3_2 _15278_ (.A(_06159_),
    .B(_06168_),
    .C(_06170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06173_));
 sky130_fd_sc_hd__a21oi_2 _15279_ (.A1(_06168_),
    .A2(_06170_),
    .B1(_06159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06174_));
 sky130_fd_sc_hd__o21bai_2 _15280_ (.A1(_06167_),
    .A2(_06169_),
    .B1_N(_06159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_2 _15281_ (.A(_06157_),
    .B(_06175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06176_));
 sky130_fd_sc_hd__a22o_2 _15282_ (.A1(_06154_),
    .A2(_06156_),
    .B1(_06173_),
    .B2(_06175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06177_));
 sky130_fd_sc_hd__o21ai_2 _15283_ (.A1(_06172_),
    .A2(_06176_),
    .B1(_06177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06178_));
 sky130_fd_sc_hd__o211ai_2 _15284_ (.A1(_06172_),
    .A2(_06176_),
    .B1(_05999_),
    .C1(_06177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06179_));
 sky130_fd_sc_hd__o21ai_2 _15285_ (.A1(_06153_),
    .A2(_06155_),
    .B1(_06175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06180_));
 sky130_fd_sc_hd__a21o_2 _15286_ (.A1(_06173_),
    .A2(_06175_),
    .B1(_06158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06181_));
 sky130_fd_sc_hd__o211ai_2 _15287_ (.A1(_06180_),
    .A2(_06172_),
    .B1(_06000_),
    .C1(_06181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06182_));
 sky130_fd_sc_hd__o22a_2 _15288_ (.A1(_06111_),
    .A2(_06112_),
    .B1(_06101_),
    .B2(_06105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06183_));
 sky130_fd_sc_hd__a2bb2o_2 _15289_ (.A1_N(_06101_),
    .A2_N(_06105_),
    .B1(_06113_),
    .B2(_06104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06184_));
 sky130_fd_sc_hd__o2bb2ai_2 _15290_ (.A1_N(_06179_),
    .A2_N(_06182_),
    .B1(_06183_),
    .B2(_06103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06185_));
 sky130_fd_sc_hd__nand3_2 _15291_ (.A(_06179_),
    .B(_06182_),
    .C(_06184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06186_));
 sky130_fd_sc_hd__nand2_2 _15292_ (.A(_06185_),
    .B(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06187_));
 sky130_fd_sc_hd__a32oi_2 _15293_ (.A1(_06122_),
    .A2(_06123_),
    .A3(_06090_),
    .B1(_06185_),
    .B2(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06188_));
 sky130_fd_sc_hd__a32o_2 _15294_ (.A1(_06122_),
    .A2(_06123_),
    .A3(_06090_),
    .B1(_06185_),
    .B2(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06189_));
 sky130_fd_sc_hd__nor2_2 _15295_ (.A(_06127_),
    .B(_06187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_2 _15296_ (.A(_06188_),
    .B(_06190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06191_));
 sky130_fd_sc_hd__and3_2 _15297_ (.A(_06110_),
    .B(\a_h[9] ),
    .C(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06192_));
 sky130_fd_sc_hd__a211o_2 _15298_ (.A1(_06009_),
    .A2(_06107_),
    .B1(_09362_),
    .C1(_09471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06193_));
 sky130_fd_sc_hd__o2111ai_2 _15299_ (.A1(_02362_),
    .A2(_05044_),
    .B1(_06119_),
    .C1(_06123_),
    .D1(_06193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06194_));
 sky130_fd_sc_hd__o2bb2ai_2 _15300_ (.A1_N(_06119_),
    .A2_N(_06123_),
    .B1(_06192_),
    .B2(_06108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06195_));
 sky130_fd_sc_hd__o2bb2ai_2 _15301_ (.A1_N(_06194_),
    .A2_N(_06195_),
    .B1(_09384_),
    .B2(_09471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06196_));
 sky130_fd_sc_hd__nand4_2 _15302_ (.A(_06194_),
    .B(_06195_),
    .C(\b_l[15] ),
    .D(\a_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_2 _15303_ (.A(_06196_),
    .B(_06197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06198_));
 sky130_fd_sc_hd__o211ai_2 _15304_ (.A1(_06188_),
    .A2(_06190_),
    .B1(_06196_),
    .C1(_06197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2_2 _15305_ (.A(_06191_),
    .B(_06198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06200_));
 sky130_fd_sc_hd__nand4_2 _15306_ (.A(_06130_),
    .B(_06135_),
    .C(_06199_),
    .D(_06200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06201_));
 sky130_fd_sc_hd__a22oi_2 _15307_ (.A1(_06130_),
    .A2(_06135_),
    .B1(_06199_),
    .B2(_06200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06202_));
 sky130_fd_sc_hd__a22o_2 _15308_ (.A1(_06130_),
    .A2(_06135_),
    .B1(_06199_),
    .B2(_06200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06203_));
 sky130_fd_sc_hd__a21bo_2 _15309_ (.A1(_06086_),
    .A2(_06083_),
    .B1_N(_06085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06204_));
 sky130_fd_sc_hd__nand3_2 _15310_ (.A(_06201_),
    .B(_06203_),
    .C(_06204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06205_));
 sky130_fd_sc_hd__a21o_2 _15311_ (.A1(_06201_),
    .A2(_06203_),
    .B1(_06204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06206_));
 sky130_fd_sc_hd__a21oi_2 _15312_ (.A1(_06201_),
    .A2(_06204_),
    .B1(_06202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06207_));
 sky130_fd_sc_hd__a21bo_2 _15313_ (.A1(_06205_),
    .A2(_06206_),
    .B1_N(_06139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06208_));
 sky130_fd_sc_hd__nand3b_2 _15314_ (.A_N(_06139_),
    .B(_06205_),
    .C(_06206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06209_));
 sky130_fd_sc_hd__inv_2 _15315_ (.A(_06209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06210_));
 sky130_fd_sc_hd__nand2_2 _15316_ (.A(_06208_),
    .B(_06209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06211_));
 sky130_fd_sc_hd__nor2_2 _15317_ (.A(_06073_),
    .B(_06146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06212_));
 sky130_fd_sc_hd__a32o_2 _15318_ (.A1(_06079_),
    .A2(_06140_),
    .A3(_06141_),
    .B1(_06071_),
    .B2(_06144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06213_));
 sky130_fd_sc_hd__a21oi_2 _15319_ (.A1(_06074_),
    .A2(_06212_),
    .B1(_06213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06214_));
 sky130_fd_sc_hd__nand2_2 _15320_ (.A(_06075_),
    .B(_06212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06215_));
 sky130_fd_sc_hd__nand2_2 _15321_ (.A(_06214_),
    .B(_06215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06216_));
 sky130_fd_sc_hd__nand3_2 _15322_ (.A(_05888_),
    .B(_05889_),
    .C(_06214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06217_));
 sky130_fd_sc_hd__nand2_2 _15323_ (.A(_06216_),
    .B(_06217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06218_));
 sky130_fd_sc_hd__a21oi_2 _15324_ (.A1(_06218_),
    .A2(_06211_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06219_));
 sky130_fd_sc_hd__o21a_2 _15325_ (.A1(_06211_),
    .A2(_06218_),
    .B1(_06219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00330_));
 sky130_fd_sc_hd__nand2_2 _15326_ (.A(_06195_),
    .B(_06197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06220_));
 sky130_fd_sc_hd__nand2_2 _15327_ (.A(\b_l[12] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06221_));
 sky130_fd_sc_hd__nand2_2 _15328_ (.A(\b_l[13] ),
    .B(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06222_));
 sky130_fd_sc_hd__nand2_2 _15329_ (.A(_06221_),
    .B(_06222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06223_));
 sky130_fd_sc_hd__nand4_2 _15330_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[12] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06224_));
 sky130_fd_sc_hd__nand4_2 _15331_ (.A(_06223_),
    .B(_06224_),
    .C(\b_l[14] ),
    .D(\a_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06225_));
 sky130_fd_sc_hd__a22o_2 _15332_ (.A1(\b_l[14] ),
    .A2(\a_h[11] ),
    .B1(_06223_),
    .B2(_06224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06226_));
 sky130_fd_sc_hd__o21ai_2 _15333_ (.A1(_06161_),
    .A2(_06165_),
    .B1(_06163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06227_));
 sky130_fd_sc_hd__nand2_2 _15334_ (.A(\b_l[11] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_2 _15335_ (.A(\b_l[11] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2_2 _15336_ (.A(_06162_),
    .B(_06228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06230_));
 sky130_fd_sc_hd__o21a_2 _15337_ (.A1(_06095_),
    .A2(_06229_),
    .B1(_06230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06231_));
 sky130_fd_sc_hd__o21ai_2 _15338_ (.A1(_06095_),
    .A2(_06229_),
    .B1(_06230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06232_));
 sky130_fd_sc_hd__o211ai_2 _15339_ (.A1(_06165_),
    .A2(_06161_),
    .B1(_06163_),
    .C1(_06232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06233_));
 sky130_fd_sc_hd__nand2_2 _15340_ (.A(_06227_),
    .B(_06231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06234_));
 sky130_fd_sc_hd__a22o_2 _15341_ (.A1(_06225_),
    .A2(_06226_),
    .B1(_06233_),
    .B2(_06234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06235_));
 sky130_fd_sc_hd__nand4_2 _15342_ (.A(_06225_),
    .B(_06226_),
    .C(_06233_),
    .D(_06234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06236_));
 sky130_fd_sc_hd__o22ai_2 _15343_ (.A1(_06167_),
    .A2(_06171_),
    .B1(_06158_),
    .B2(_06174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06237_));
 sky130_fd_sc_hd__nand3_2 _15344_ (.A(_06237_),
    .B(_06236_),
    .C(_06235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06238_));
 sky130_fd_sc_hd__a221o_2 _15345_ (.A1(_06157_),
    .A2(_06175_),
    .B1(_06235_),
    .B2(_06236_),
    .C1(_06172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06239_));
 sky130_fd_sc_hd__and2_2 _15346_ (.A(_06238_),
    .B(_06239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06240_));
 sky130_fd_sc_hd__nor2_2 _15347_ (.A(_09384_),
    .B(_09482_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06241_));
 sky130_fd_sc_hd__o31a_2 _15348_ (.A1(_09362_),
    .A2(_09482_),
    .A3(_06149_),
    .B1(_06152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06242_));
 sky130_fd_sc_hd__a2bb2oi_2 _15349_ (.A1_N(_06151_),
    .A2_N(_06155_),
    .B1(_06179_),
    .B2(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06243_));
 sky130_fd_sc_hd__a21o_2 _15350_ (.A1(_06179_),
    .A2(_06186_),
    .B1(_06242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06244_));
 sky130_fd_sc_hd__o211a_2 _15351_ (.A1(_06000_),
    .A2(_06178_),
    .B1(_06242_),
    .C1(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06245_));
 sky130_fd_sc_hd__o211ai_2 _15352_ (.A1(_06000_),
    .A2(_06178_),
    .B1(_06242_),
    .C1(_06186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06246_));
 sky130_fd_sc_hd__o22ai_2 _15353_ (.A1(_09384_),
    .A2(_09482_),
    .B1(_06243_),
    .B2(_06245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06247_));
 sky130_fd_sc_hd__nand3_2 _15354_ (.A(_06244_),
    .B(_06246_),
    .C(_06241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06248_));
 sky130_fd_sc_hd__a21oi_2 _15355_ (.A1(_06247_),
    .A2(_06248_),
    .B1(_06240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06249_));
 sky130_fd_sc_hd__and3_2 _15356_ (.A(_06247_),
    .B(_06248_),
    .C(_06240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06250_));
 sky130_fd_sc_hd__nand3_2 _15357_ (.A(_06247_),
    .B(_06248_),
    .C(_06240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06251_));
 sky130_fd_sc_hd__a31o_2 _15358_ (.A1(_06189_),
    .A2(_06196_),
    .A3(_06197_),
    .B1(_06190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06252_));
 sky130_fd_sc_hd__o21bai_2 _15359_ (.A1(_06249_),
    .A2(_06250_),
    .B1_N(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06253_));
 sky130_fd_sc_hd__nand3b_2 _15360_ (.A_N(_06249_),
    .B(_06251_),
    .C(_06252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06254_));
 sky130_fd_sc_hd__a21oi_2 _15361_ (.A1(_06253_),
    .A2(_06254_),
    .B1(_06220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06255_));
 sky130_fd_sc_hd__and3_2 _15362_ (.A(_06220_),
    .B(_06253_),
    .C(_06254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06256_));
 sky130_fd_sc_hd__nand3_2 _15363_ (.A(_06220_),
    .B(_06253_),
    .C(_06254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06257_));
 sky130_fd_sc_hd__o21ai_2 _15364_ (.A1(_06255_),
    .A2(_06256_),
    .B1(_06207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06258_));
 sky130_fd_sc_hd__nor2_2 _15365_ (.A(_06207_),
    .B(_06255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06259_));
 sky130_fd_sc_hd__nand2_2 _15366_ (.A(_06259_),
    .B(_06257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_2 _15367_ (.A(_06258_),
    .B(_06260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06261_));
 sky130_fd_sc_hd__a31oi_2 _15368_ (.A1(_06208_),
    .A2(_06216_),
    .A3(_06217_),
    .B1(_06210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06262_));
 sky130_fd_sc_hd__o21ai_2 _15369_ (.A1(_06261_),
    .A2(_06262_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06263_));
 sky130_fd_sc_hd__a21oi_2 _15370_ (.A1(_06261_),
    .A2(_06262_),
    .B1(_06263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_2 _15371_ (.A(\b_l[13] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06264_));
 sky130_fd_sc_hd__nand2_2 _15372_ (.A(\b_l[13] ),
    .B(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06265_));
 sky130_fd_sc_hd__nand2_2 _15373_ (.A(\b_l[12] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06266_));
 sky130_fd_sc_hd__nand4_2 _15374_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[13] ),
    .D(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06267_));
 sky130_fd_sc_hd__nand2_2 _15375_ (.A(_06265_),
    .B(_06266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06268_));
 sky130_fd_sc_hd__o2111ai_2 _15376_ (.A1(_06221_),
    .A2(_06264_),
    .B1(\b_l[14] ),
    .C1(\a_h[12] ),
    .D1(_06268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06269_));
 sky130_fd_sc_hd__a22o_2 _15377_ (.A1(\b_l[14] ),
    .A2(\a_h[12] ),
    .B1(_06267_),
    .B2(_06268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06270_));
 sky130_fd_sc_hd__a32o_2 _15378_ (.A1(\b_l[11] ),
    .A2(_06095_),
    .A3(\a_h[15] ),
    .B1(_06270_),
    .B2(_06269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06271_));
 sky130_fd_sc_hd__nand4b_2 _15379_ (.A_N(_06229_),
    .B(_06269_),
    .C(_06270_),
    .D(_06095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06272_));
 sky130_fd_sc_hd__a22o_2 _15380_ (.A1(_06231_),
    .A2(_06227_),
    .B1(_06226_),
    .B2(_06225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06273_));
 sky130_fd_sc_hd__o21a_2 _15381_ (.A1(_06227_),
    .A2(_06231_),
    .B1(_06273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06274_));
 sky130_fd_sc_hd__nand4_2 _15382_ (.A(_06233_),
    .B(_06271_),
    .C(_06272_),
    .D(_06273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06275_));
 sky130_fd_sc_hd__a22o_2 _15383_ (.A1(_06271_),
    .A2(_06272_),
    .B1(_06273_),
    .B2(_06233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06276_));
 sky130_fd_sc_hd__nand2_2 _15384_ (.A(_06275_),
    .B(_06276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06277_));
 sky130_fd_sc_hd__o31a_2 _15385_ (.A1(_09504_),
    .A2(_09515_),
    .A3(_05044_),
    .B1(_06225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06278_));
 sky130_fd_sc_hd__o21ai_2 _15386_ (.A1(_06221_),
    .A2(_06222_),
    .B1(_06225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06279_));
 sky130_fd_sc_hd__o311a_2 _15387_ (.A1(_09504_),
    .A2(_09515_),
    .A3(_05044_),
    .B1(_06225_),
    .C1(_06238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06280_));
 sky130_fd_sc_hd__nand2_2 _15388_ (.A(_06238_),
    .B(_06278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06281_));
 sky130_fd_sc_hd__nand4_2 _15389_ (.A(_06237_),
    .B(_06279_),
    .C(_06235_),
    .D(_06236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06282_));
 sky130_fd_sc_hd__a22oi_2 _15390_ (.A1(\b_l[15] ),
    .A2(\a_h[11] ),
    .B1(_06281_),
    .B2(_06282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06283_));
 sky130_fd_sc_hd__nand3_2 _15391_ (.A(_06282_),
    .B(\a_h[11] ),
    .C(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06284_));
 sky130_fd_sc_hd__a21oi_2 _15392_ (.A1(_06238_),
    .A2(_06278_),
    .B1(_06284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06285_));
 sky130_fd_sc_hd__o21ai_2 _15393_ (.A1(_06283_),
    .A2(_06285_),
    .B1(_06277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06286_));
 sky130_fd_sc_hd__a41o_2 _15394_ (.A1(\b_l[15] ),
    .A2(_06281_),
    .A3(_06282_),
    .A4(\a_h[11] ),
    .B1(_06277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06287_));
 sky130_fd_sc_hd__nor2_2 _15395_ (.A(_06283_),
    .B(_06287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06288_));
 sky130_fd_sc_hd__o21a_2 _15396_ (.A1(_06283_),
    .A2(_06287_),
    .B1(_06286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06289_));
 sky130_fd_sc_hd__o21ai_2 _15397_ (.A1(_06283_),
    .A2(_06287_),
    .B1(_06286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06290_));
 sky130_fd_sc_hd__a31oi_2 _15398_ (.A1(_06247_),
    .A2(_06248_),
    .A3(_06240_),
    .B1(_06289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2_2 _15399_ (.A(_06251_),
    .B(_06290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06292_));
 sky130_fd_sc_hd__nand4_2 _15400_ (.A(_06247_),
    .B(_06289_),
    .C(_06248_),
    .D(_06240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06293_));
 sky130_fd_sc_hd__nand2_2 _15401_ (.A(_06292_),
    .B(_06293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06294_));
 sky130_fd_sc_hd__a31o_2 _15402_ (.A1(_06246_),
    .A2(\a_h[10] ),
    .A3(\b_l[15] ),
    .B1(_06243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06295_));
 sky130_fd_sc_hd__o21bai_2 _15403_ (.A1(_06251_),
    .A2(_06290_),
    .B1_N(_06295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06296_));
 sky130_fd_sc_hd__o2bb2ai_2 _15404_ (.A1_N(_06295_),
    .A2_N(_06294_),
    .B1(_06291_),
    .B2(_06296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06297_));
 sky130_fd_sc_hd__a21boi_2 _15405_ (.A1(_06254_),
    .A2(_06257_),
    .B1_N(_06297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06298_));
 sky130_fd_sc_hd__a21bo_2 _15406_ (.A1(_06254_),
    .A2(_06257_),
    .B1_N(_06297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06299_));
 sky130_fd_sc_hd__nand3b_2 _15407_ (.A_N(_06297_),
    .B(_06257_),
    .C(_06254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_2 _15408_ (.A(_06299_),
    .B(_06300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06301_));
 sky130_fd_sc_hd__and4_2 _15409_ (.A(_06208_),
    .B(_06209_),
    .C(_06258_),
    .D(_06260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06302_));
 sky130_fd_sc_hd__a21boi_2 _15410_ (.A1(_06214_),
    .A2(_06215_),
    .B1_N(_06302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06303_));
 sky130_fd_sc_hd__nand2_2 _15411_ (.A(_06217_),
    .B(_06303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06304_));
 sky130_fd_sc_hd__a22oi_2 _15412_ (.A1(_06257_),
    .A2(_06259_),
    .B1(_06210_),
    .B2(_06258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06305_));
 sky130_fd_sc_hd__a21boi_2 _15413_ (.A1(_06217_),
    .A2(_06303_),
    .B1_N(_06305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06306_));
 sky130_fd_sc_hd__and3_2 _15414_ (.A(_06301_),
    .B(_06304_),
    .C(_06305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06307_));
 sky130_fd_sc_hd__a21oi_2 _15415_ (.A1(_06304_),
    .A2(_06305_),
    .B1(_06301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06308_));
 sky130_fd_sc_hd__nor3_2 _15416_ (.A(rst),
    .B(_06307_),
    .C(_06308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00332_));
 sky130_fd_sc_hd__o21ai_2 _15417_ (.A1(_06250_),
    .A2(_06289_),
    .B1(_06296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06309_));
 sky130_fd_sc_hd__a22o_2 _15418_ (.A1(\b_l[13] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06310_));
 sky130_fd_sc_hd__nand4_2 _15419_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06311_));
 sky130_fd_sc_hd__and4_2 _15420_ (.A(_06310_),
    .B(_06311_),
    .C(\b_l[14] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06312_));
 sky130_fd_sc_hd__o2bb2a_2 _15421_ (.A1_N(_06310_),
    .A2_N(_06311_),
    .B1(_09362_),
    .B2(_09515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06313_));
 sky130_fd_sc_hd__nor2_2 _15422_ (.A(_06312_),
    .B(_06313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06314_));
 sky130_fd_sc_hd__o21ai_2 _15423_ (.A1(_06095_),
    .A2(_06229_),
    .B1(_06272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06315_));
 sky130_fd_sc_hd__xor2_2 _15424_ (.A(_06314_),
    .B(_06315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06316_));
 sky130_fd_sc_hd__o31a_2 _15425_ (.A1(_09351_),
    .A2(_09515_),
    .A3(_06266_),
    .B1(_06269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06317_));
 sky130_fd_sc_hd__o21ai_2 _15426_ (.A1(_06265_),
    .A2(_06266_),
    .B1(_06269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06318_));
 sky130_fd_sc_hd__and4_2 _15427_ (.A(_06274_),
    .B(_06318_),
    .C(_06271_),
    .D(_06272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06319_));
 sky130_fd_sc_hd__nand4_2 _15428_ (.A(_06274_),
    .B(_06318_),
    .C(_06271_),
    .D(_06272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_2 _15429_ (.A(_06275_),
    .B(_06317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06321_));
 sky130_fd_sc_hd__nand4_2 _15430_ (.A(_06320_),
    .B(_06321_),
    .C(\b_l[15] ),
    .D(\a_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06322_));
 sky130_fd_sc_hd__a22o_2 _15431_ (.A1(\b_l[15] ),
    .A2(\a_h[12] ),
    .B1(_06320_),
    .B2(_06321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06323_));
 sky130_fd_sc_hd__nand3_2 _15432_ (.A(_06323_),
    .B(_06316_),
    .C(_06322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06324_));
 sky130_fd_sc_hd__a21o_2 _15433_ (.A1(_06322_),
    .A2(_06323_),
    .B1(_06316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06325_));
 sky130_fd_sc_hd__a2bb2o_2 _15434_ (.A1_N(_06283_),
    .A2_N(_06287_),
    .B1(_06324_),
    .B2(_06325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06326_));
 sky130_fd_sc_hd__nand3_2 _15435_ (.A(_06325_),
    .B(_06288_),
    .C(_06324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06327_));
 sky130_fd_sc_hd__o31ai_2 _15436_ (.A1(_09384_),
    .A2(_09493_),
    .A3(_06280_),
    .B1(_06282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06328_));
 sky130_fd_sc_hd__a21o_2 _15437_ (.A1(_06326_),
    .A2(_06327_),
    .B1(_06328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06329_));
 sky130_fd_sc_hd__nand3_2 _15438_ (.A(_06326_),
    .B(_06327_),
    .C(_06328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06330_));
 sky130_fd_sc_hd__and2_2 _15439_ (.A(_06329_),
    .B(_06330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06331_));
 sky130_fd_sc_hd__a22o_2 _15440_ (.A1(_06292_),
    .A2(_06296_),
    .B1(_06329_),
    .B2(_06330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06332_));
 sky130_fd_sc_hd__and3_2 _15441_ (.A(_06292_),
    .B(_06296_),
    .C(_06331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06333_));
 sky130_fd_sc_hd__xnor2_2 _15442_ (.A(_06309_),
    .B(_06331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06334_));
 sky130_fd_sc_hd__inv_2 _15443_ (.A(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06335_));
 sky130_fd_sc_hd__o21ai_2 _15444_ (.A1(_06301_),
    .A2(_06306_),
    .B1(_06335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06336_));
 sky130_fd_sc_hd__o21ai_2 _15445_ (.A1(_06298_),
    .A2(_06308_),
    .B1(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06337_));
 sky130_fd_sc_hd__o211a_2 _15446_ (.A1(_06336_),
    .A2(_06298_),
    .B1(_09690_),
    .C1(_06337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00333_));
 sky130_fd_sc_hd__and2b_2 _15447_ (.A_N(_06301_),
    .B(_06334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06338_));
 sky130_fd_sc_hd__nand2_2 _15448_ (.A(_06302_),
    .B(_06338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06339_));
 sky130_fd_sc_hd__a21oi_2 _15449_ (.A1(_06214_),
    .A2(_06215_),
    .B1(_06339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06340_));
 sky130_fd_sc_hd__nand2_2 _15450_ (.A(_06217_),
    .B(_06340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06341_));
 sky130_fd_sc_hd__o21ai_2 _15451_ (.A1(_06298_),
    .A2(_06333_),
    .B1(_06332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06342_));
 sky130_fd_sc_hd__o31a_2 _15452_ (.A1(_06301_),
    .A2(_06305_),
    .A3(_06335_),
    .B1(_06342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06343_));
 sky130_fd_sc_hd__o31ai_2 _15453_ (.A1(_06301_),
    .A2(_06305_),
    .A3(_06335_),
    .B1(_06342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06344_));
 sky130_fd_sc_hd__a21oi_2 _15454_ (.A1(_06217_),
    .A2(_06340_),
    .B1(_06344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06345_));
 sky130_fd_sc_hd__a21boi_2 _15455_ (.A1(_06326_),
    .A2(_06328_),
    .B1_N(_06327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06346_));
 sky130_fd_sc_hd__a22oi_2 _15456_ (.A1(\b_l[14] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06347_));
 sky130_fd_sc_hd__and4_2 _15457_ (.A(\b_l[13] ),
    .B(\b_l[14] ),
    .C(\a_h[14] ),
    .D(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06348_));
 sky130_fd_sc_hd__a31o_2 _15458_ (.A1(\a_h[14] ),
    .A2(\a_h[15] ),
    .A3(_05043_),
    .B1(_06312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06349_));
 sky130_fd_sc_hd__a21oi_2 _15459_ (.A1(_06315_),
    .A2(_06314_),
    .B1(_06349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06350_));
 sky130_fd_sc_hd__nand3_2 _15460_ (.A(_06315_),
    .B(_06349_),
    .C(_06314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06351_));
 sky130_fd_sc_hd__inv_2 _15461_ (.A(_06351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06352_));
 sky130_fd_sc_hd__and4b_2 _15462_ (.A_N(_06350_),
    .B(_06351_),
    .C(\b_l[15] ),
    .D(\a_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06353_));
 sky130_fd_sc_hd__o22a_2 _15463_ (.A1(_09384_),
    .A2(_09515_),
    .B1(_06350_),
    .B2(_06352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06354_));
 sky130_fd_sc_hd__nor4_2 _15464_ (.A(_06347_),
    .B(_06348_),
    .C(_06353_),
    .D(_06354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06355_));
 sky130_fd_sc_hd__o22ai_2 _15465_ (.A1(_06347_),
    .A2(_06348_),
    .B1(_06353_),
    .B2(_06354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06356_));
 sky130_fd_sc_hd__inv_2 _15466_ (.A(_06356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06357_));
 sky130_fd_sc_hd__o21a_2 _15467_ (.A1(_06355_),
    .A2(_06357_),
    .B1(_06324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06358_));
 sky130_fd_sc_hd__nor3_2 _15468_ (.A(_06324_),
    .B(_06355_),
    .C(_06357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06359_));
 sky130_fd_sc_hd__a31o_2 _15469_ (.A1(\b_l[15] ),
    .A2(\a_h[12] ),
    .A3(_06321_),
    .B1(_06319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06360_));
 sky130_fd_sc_hd__o21ai_2 _15470_ (.A1(_06358_),
    .A2(_06359_),
    .B1(_06360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06361_));
 sky130_fd_sc_hd__or3_2 _15471_ (.A(_06358_),
    .B(_06359_),
    .C(_06360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06362_));
 sky130_fd_sc_hd__nand2_2 _15472_ (.A(_06361_),
    .B(_06362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06363_));
 sky130_fd_sc_hd__and2b_2 _15473_ (.A_N(_06346_),
    .B(_06363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06364_));
 sky130_fd_sc_hd__xor2_2 _15474_ (.A(_06346_),
    .B(_06363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06365_));
 sky130_fd_sc_hd__a21oi_2 _15475_ (.A1(_06341_),
    .A2(_06343_),
    .B1(_06365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06366_));
 sky130_fd_sc_hd__o21ai_2 _15476_ (.A1(_06365_),
    .A2(_06345_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06367_));
 sky130_fd_sc_hd__a21oi_2 _15477_ (.A1(_06345_),
    .A2(_06365_),
    .B1(_06367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00334_));
 sky130_fd_sc_hd__a31o_2 _15478_ (.A1(_06314_),
    .A2(_06315_),
    .A3(_06349_),
    .B1(_06353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06368_));
 sky130_fd_sc_hd__nand2_2 _15479_ (.A(\b_l[14] ),
    .B(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06369_));
 sky130_fd_sc_hd__nand2_2 _15480_ (.A(\b_l[15] ),
    .B(\a_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06370_));
 sky130_fd_sc_hd__o22a_2 _15481_ (.A1(\b_l[15] ),
    .A2(_06264_),
    .B1(_06370_),
    .B2(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06371_));
 sky130_fd_sc_hd__or3b_2 _15482_ (.A(_09362_),
    .B(_06371_),
    .C_N(\a_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06372_));
 sky130_fd_sc_hd__a22o_2 _15483_ (.A1(\b_l[15] ),
    .A2(\a_h[14] ),
    .B1(\a_h[15] ),
    .B2(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06373_));
 sky130_fd_sc_hd__a21o_2 _15484_ (.A1(_06372_),
    .A2(_06373_),
    .B1(_06355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06374_));
 sky130_fd_sc_hd__inv_2 _15485_ (.A(_06374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06375_));
 sky130_fd_sc_hd__and3_2 _15486_ (.A(_06355_),
    .B(_06372_),
    .C(_06373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06376_));
 sky130_fd_sc_hd__o22a_2 _15487_ (.A1(_06352_),
    .A2(_06353_),
    .B1(_06375_),
    .B2(_06376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06377_));
 sky130_fd_sc_hd__o21ai_2 _15488_ (.A1(_06375_),
    .A2(_06376_),
    .B1(_06368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06378_));
 sky130_fd_sc_hd__or3_2 _15489_ (.A(_06376_),
    .B(_06368_),
    .C(_06375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06379_));
 sky130_fd_sc_hd__nand2b_2 _15490_ (.A_N(_06358_),
    .B(_06360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06380_));
 sky130_fd_sc_hd__inv_2 _15491_ (.A(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06381_));
 sky130_fd_sc_hd__o2bb2a_2 _15492_ (.A1_N(_06378_),
    .A2_N(_06379_),
    .B1(_06381_),
    .B2(_06359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06382_));
 sky130_fd_sc_hd__or4bb_2 _15493_ (.A(_06359_),
    .B(_06377_),
    .C_N(_06379_),
    .D_N(_06380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06383_));
 sky130_fd_sc_hd__nand2b_2 _15494_ (.A_N(_06382_),
    .B(_06383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06384_));
 sky130_fd_sc_hd__o21ai_2 _15495_ (.A1(_06365_),
    .A2(_06345_),
    .B1(_06384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06385_));
 sky130_fd_sc_hd__o21bai_2 _15496_ (.A1(_06364_),
    .A2(_06366_),
    .B1_N(_06384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06386_));
 sky130_fd_sc_hd__o211a_2 _15497_ (.A1(_06385_),
    .A2(_06364_),
    .B1(_09690_),
    .C1(_06386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00335_));
 sky130_fd_sc_hd__o2bb2a_2 _15498_ (.A1_N(\b_l[15] ),
    .A2_N(\a_h[15] ),
    .B1(_06369_),
    .B2(_06371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06387_));
 sky130_fd_sc_hd__a41o_2 _15499_ (.A1(\b_l[14] ),
    .A2(\b_l[15] ),
    .A3(\a_h[14] ),
    .A4(\a_h[15] ),
    .B1(_06387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06388_));
 sky130_fd_sc_hd__a21oi_2 _15500_ (.A1(_06368_),
    .A2(_06374_),
    .B1(_06376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06389_));
 sky130_fd_sc_hd__xor2_2 _15501_ (.A(_06388_),
    .B(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06390_));
 sky130_fd_sc_hd__inv_2 _15502_ (.A(_06390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06391_));
 sky130_fd_sc_hd__o21a_2 _15503_ (.A1(_06364_),
    .A2(_06382_),
    .B1(_06383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06392_));
 sky130_fd_sc_hd__inv_2 _15504_ (.A(_06392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06393_));
 sky130_fd_sc_hd__or2_2 _15505_ (.A(_06365_),
    .B(_06384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06394_));
 sky130_fd_sc_hd__a21oi_2 _15506_ (.A1(_06341_),
    .A2(_06343_),
    .B1(_06394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06395_));
 sky130_fd_sc_hd__o211ai_2 _15507_ (.A1(_06394_),
    .A2(_06345_),
    .B1(_06391_),
    .C1(_06393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06396_));
 sky130_fd_sc_hd__o21a_2 _15508_ (.A1(_06392_),
    .A2(_06395_),
    .B1(_06390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06397_));
 sky130_fd_sc_hd__o21ai_2 _15509_ (.A1(_06392_),
    .A2(_06395_),
    .B1(_06390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06398_));
 sky130_fd_sc_hd__nand2_2 _15510_ (.A(_09690_),
    .B(_06396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06399_));
 sky130_fd_sc_hd__nor2_2 _15511_ (.A(_06397_),
    .B(_06399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00336_));
 sky130_fd_sc_hd__o22a_2 _15512_ (.A1(_06369_),
    .A2(_06370_),
    .B1(_06387_),
    .B2(_06389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06400_));
 sky130_fd_sc_hd__a21oi_2 _15513_ (.A1(_06398_),
    .A2(_06400_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00337_));
 sky130_fd_sc_hd__and3_2 _15514_ (.A(_09690_),
    .B(\b_h[0] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00338_));
 sky130_fd_sc_hd__and2_2 _15515_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06401_));
 sky130_fd_sc_hd__nand2_2 _15516_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06402_));
 sky130_fd_sc_hd__o2bb2a_2 _15517_ (.A1_N(\a_l[1] ),
    .A2_N(\b_h[0] ),
    .B1(_09581_),
    .B2(_09166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06403_));
 sky130_fd_sc_hd__a311oi_2 _15518_ (.A1(\b_h[0] ),
    .A2(\b_h[1] ),
    .A3(_06401_),
    .B1(_06403_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00339_));
 sky130_fd_sc_hd__or3_2 _15519_ (.A(_09581_),
    .B(_09592_),
    .C(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06404_));
 sky130_fd_sc_hd__a22o_2 _15520_ (.A1(\a_l[1] ),
    .A2(\b_h[1] ),
    .B1(\b_h[2] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06405_));
 sky130_fd_sc_hd__nand4_2 _15521_ (.A(_06404_),
    .B(_06405_),
    .C(\a_l[2] ),
    .D(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06406_));
 sky130_fd_sc_hd__a22o_2 _15522_ (.A1(\a_l[2] ),
    .A2(\b_h[0] ),
    .B1(_06404_),
    .B2(_06405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06407_));
 sky130_fd_sc_hd__nand2_2 _15523_ (.A(_06406_),
    .B(_06407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06408_));
 sky130_fd_sc_hd__o31a_2 _15524_ (.A1(_09526_),
    .A2(_09581_),
    .A3(_06402_),
    .B1(_06408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06409_));
 sky130_fd_sc_hd__and4_2 _15525_ (.A(_06407_),
    .B(_01856_),
    .C(_06406_),
    .D(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06410_));
 sky130_fd_sc_hd__nor3_2 _15526_ (.A(rst),
    .B(_06409_),
    .C(_06410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_2 _15527_ (.A(\a_l[3] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_2 _15528_ (.A(\a_l[2] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06412_));
 sky130_fd_sc_hd__nand2_2 _15529_ (.A(\a_l[1] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06413_));
 sky130_fd_sc_hd__nand4_2 _15530_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06414_));
 sky130_fd_sc_hd__a22oi_2 _15531_ (.A1(\a_l[1] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06415_));
 sky130_fd_sc_hd__a22o_2 _15532_ (.A1(\a_l[1] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06416_));
 sky130_fd_sc_hd__o211a_2 _15533_ (.A1(_09144_),
    .A2(_09581_),
    .B1(_06414_),
    .C1(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06417_));
 sky130_fd_sc_hd__o211ai_2 _15534_ (.A1(_09144_),
    .A2(_09581_),
    .B1(_06414_),
    .C1(_06416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06418_));
 sky130_fd_sc_hd__a21oi_2 _15535_ (.A1(_06414_),
    .A2(_06416_),
    .B1(_06412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06419_));
 sky130_fd_sc_hd__a21o_2 _15536_ (.A1(_06414_),
    .A2(_06416_),
    .B1(_06412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06420_));
 sky130_fd_sc_hd__o21bai_2 _15537_ (.A1(_06417_),
    .A2(_06419_),
    .B1_N(_06404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06421_));
 sky130_fd_sc_hd__nand3_2 _15538_ (.A(_06404_),
    .B(_06418_),
    .C(_06420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06422_));
 sky130_fd_sc_hd__o211ai_2 _15539_ (.A1(_09188_),
    .A2(_09526_),
    .B1(_06421_),
    .C1(_06422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06423_));
 sky130_fd_sc_hd__a21o_2 _15540_ (.A1(_06421_),
    .A2(_06422_),
    .B1(_06411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06424_));
 sky130_fd_sc_hd__nand3_2 _15541_ (.A(_06406_),
    .B(_06423_),
    .C(_06424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06425_));
 sky130_fd_sc_hd__or4b_2 _15542_ (.A(_01857_),
    .B(_06402_),
    .C(_06408_),
    .D_N(_06425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06426_));
 sky130_fd_sc_hd__a21oi_2 _15543_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06427_));
 sky130_fd_sc_hd__a21o_2 _15544_ (.A1(_06423_),
    .A2(_06424_),
    .B1(_06406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06428_));
 sky130_fd_sc_hd__a21o_2 _15545_ (.A1(_06425_),
    .A2(_06428_),
    .B1(_06410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06429_));
 sky130_fd_sc_hd__and3_2 _15546_ (.A(_09690_),
    .B(_06426_),
    .C(_06429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00341_));
 sky130_fd_sc_hd__a32o_2 _15547_ (.A1(_06404_),
    .A2(_06418_),
    .A3(_06420_),
    .B1(_06421_),
    .B2(_06411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06430_));
 sky130_fd_sc_hd__nand2_2 _15548_ (.A(\a_l[4] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2_2 _15549_ (.A(\a_l[0] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06432_));
 sky130_fd_sc_hd__and4_2 _15550_ (.A(\a_l[0] ),
    .B(\a_l[4] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06433_));
 sky130_fd_sc_hd__o21a_2 _15551_ (.A1(_09199_),
    .A2(_09526_),
    .B1(_06432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06434_));
 sky130_fd_sc_hd__or2_2 _15552_ (.A(_06433_),
    .B(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06435_));
 sky130_fd_sc_hd__a21oi_2 _15553_ (.A1(_06412_),
    .A2(_06414_),
    .B1(_06415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06436_));
 sky130_fd_sc_hd__and2_2 _15554_ (.A(\a_l[3] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06437_));
 sky130_fd_sc_hd__nand2_2 _15555_ (.A(\a_l[2] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06438_));
 sky130_fd_sc_hd__nand2_2 _15556_ (.A(_06413_),
    .B(_06438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06439_));
 sky130_fd_sc_hd__nand2_2 _15557_ (.A(\b_h[2] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_2 _15558_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06441_));
 sky130_fd_sc_hd__nand4_2 _15559_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06442_));
 sky130_fd_sc_hd__and3_2 _15560_ (.A(_06439_),
    .B(_06442_),
    .C(_06437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06443_));
 sky130_fd_sc_hd__o2111ai_2 _15561_ (.A1(_06440_),
    .A2(_06441_),
    .B1(\a_l[3] ),
    .C1(\b_h[1] ),
    .D1(_06439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06444_));
 sky130_fd_sc_hd__a21oi_2 _15562_ (.A1(_06439_),
    .A2(_06442_),
    .B1(_06437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06445_));
 sky130_fd_sc_hd__a21o_2 _15563_ (.A1(_06439_),
    .A2(_06442_),
    .B1(_06437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06446_));
 sky130_fd_sc_hd__nand3_2 _15564_ (.A(_06446_),
    .B(_06436_),
    .C(_06444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06447_));
 sky130_fd_sc_hd__a21oi_2 _15565_ (.A1(_06444_),
    .A2(_06446_),
    .B1(_06436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06448_));
 sky130_fd_sc_hd__o21bai_2 _15566_ (.A1(_06443_),
    .A2(_06445_),
    .B1_N(_06436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06449_));
 sky130_fd_sc_hd__and3_2 _15567_ (.A(_06435_),
    .B(_06447_),
    .C(_06449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06450_));
 sky130_fd_sc_hd__o211ai_2 _15568_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06447_),
    .C1(_06449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06451_));
 sky130_fd_sc_hd__a21oi_2 _15569_ (.A1(_06447_),
    .A2(_06449_),
    .B1(_06435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06452_));
 sky130_fd_sc_hd__a211o_2 _15570_ (.A1(_06447_),
    .A2(_06449_),
    .B1(_06433_),
    .C1(_06434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06453_));
 sky130_fd_sc_hd__nand3_2 _15571_ (.A(_06430_),
    .B(_06451_),
    .C(_06453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06454_));
 sky130_fd_sc_hd__o21bai_2 _15572_ (.A1(_06450_),
    .A2(_06452_),
    .B1_N(_06430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2_2 _15573_ (.A(_06454_),
    .B(_06455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06456_));
 sky130_fd_sc_hd__and3_2 _15574_ (.A(_06426_),
    .B(_06428_),
    .C(_06456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06457_));
 sky130_fd_sc_hd__and4_2 _15575_ (.A(_06425_),
    .B(_06454_),
    .C(_06455_),
    .D(_06410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06458_));
 sky130_fd_sc_hd__nand2_2 _15576_ (.A(_06454_),
    .B(_06427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06459_));
 sky130_fd_sc_hd__and4_2 _15577_ (.A(_06425_),
    .B(_06454_),
    .C(_06455_),
    .D(_06410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06460_));
 sky130_fd_sc_hd__nor4b_2 _15578_ (.A(rst),
    .B(_06457_),
    .C(_06458_),
    .D_N(_06459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00342_));
 sky130_fd_sc_hd__o21a_2 _15579_ (.A1(_06433_),
    .A2(_06434_),
    .B1(_06447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06461_));
 sky130_fd_sc_hd__o21ai_2 _15580_ (.A1(_06435_),
    .A2(_06448_),
    .B1(_06447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_2 _15581_ (.A(\a_l[0] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_2 _15582_ (.A(\a_l[1] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06464_));
 sky130_fd_sc_hd__nand2_2 _15583_ (.A(\a_l[5] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06465_));
 sky130_fd_sc_hd__nand2_2 _15584_ (.A(_06464_),
    .B(_06465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_2 _15585_ (.A(\a_l[5] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06467_));
 sky130_fd_sc_hd__and4_2 _15586_ (.A(\a_l[1] ),
    .B(\a_l[5] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06468_));
 sky130_fd_sc_hd__nand4_2 _15587_ (.A(\a_l[1] ),
    .B(\a_l[5] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06469_));
 sky130_fd_sc_hd__a21o_2 _15588_ (.A1(_06466_),
    .A2(_06469_),
    .B1(_06463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06470_));
 sky130_fd_sc_hd__o211ai_2 _15589_ (.A1(_09166_),
    .A2(_09602_),
    .B1(_06466_),
    .C1(_06469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06471_));
 sky130_fd_sc_hd__nand2_2 _15590_ (.A(_06470_),
    .B(_06471_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06472_));
 sky130_fd_sc_hd__a21boi_2 _15591_ (.A1(_06439_),
    .A2(_06437_),
    .B1_N(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06473_));
 sky130_fd_sc_hd__a21bo_2 _15592_ (.A1(_06439_),
    .A2(_06437_),
    .B1_N(_06442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06474_));
 sky130_fd_sc_hd__nand2_2 _15593_ (.A(\a_l[4] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_2 _15594_ (.A(\a_l[2] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06476_));
 sky130_fd_sc_hd__nand2_2 _15595_ (.A(\a_l[3] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06477_));
 sky130_fd_sc_hd__a22oi_2 _15596_ (.A1(\a_l[3] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06478_));
 sky130_fd_sc_hd__nand2_2 _15597_ (.A(_06476_),
    .B(_06477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06479_));
 sky130_fd_sc_hd__nand2_2 _15598_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06480_));
 sky130_fd_sc_hd__nand4_2 _15599_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06481_));
 sky130_fd_sc_hd__o2bb2a_2 _15600_ (.A1_N(_06479_),
    .A2_N(_06481_),
    .B1(_09199_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06482_));
 sky130_fd_sc_hd__o2bb2ai_2 _15601_ (.A1_N(_06479_),
    .A2_N(_06481_),
    .B1(_09199_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06483_));
 sky130_fd_sc_hd__o2111ai_2 _15602_ (.A1(_06440_),
    .A2(_06480_),
    .B1(\a_l[4] ),
    .C1(\b_h[1] ),
    .D1(_06479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06484_));
 sky130_fd_sc_hd__a21o_2 _15603_ (.A1(_06479_),
    .A2(_06481_),
    .B1(_06475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_2 _15604_ (.A(_06475_),
    .B(_06481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06486_));
 sky130_fd_sc_hd__o221ai_2 _15605_ (.A1(_09199_),
    .A2(_09581_),
    .B1(_06440_),
    .B2(_06480_),
    .C1(_06479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06487_));
 sky130_fd_sc_hd__nand2_2 _15606_ (.A(_06474_),
    .B(_06484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06488_));
 sky130_fd_sc_hd__nand3_2 _15607_ (.A(_06474_),
    .B(_06483_),
    .C(_06484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06489_));
 sky130_fd_sc_hd__nand3_2 _15608_ (.A(_06485_),
    .B(_06487_),
    .C(_06473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06490_));
 sky130_fd_sc_hd__nand4_2 _15609_ (.A(_06470_),
    .B(_06471_),
    .C(_06489_),
    .D(_06490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06491_));
 sky130_fd_sc_hd__a22o_2 _15610_ (.A1(_06470_),
    .A2(_06471_),
    .B1(_06489_),
    .B2(_06490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06492_));
 sky130_fd_sc_hd__o211ai_2 _15611_ (.A1(_06448_),
    .A2(_06461_),
    .B1(_06491_),
    .C1(_06492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06493_));
 sky130_fd_sc_hd__o211ai_2 _15612_ (.A1(_06482_),
    .A2(_06488_),
    .B1(_06490_),
    .C1(_06472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06494_));
 sky130_fd_sc_hd__a21o_2 _15613_ (.A1(_06489_),
    .A2(_06490_),
    .B1(_06472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06495_));
 sky130_fd_sc_hd__nand3_2 _15614_ (.A(_06462_),
    .B(_06494_),
    .C(_06495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06496_));
 sky130_fd_sc_hd__nand3_2 _15615_ (.A(_06496_),
    .B(_06433_),
    .C(_06493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06497_));
 sky130_fd_sc_hd__o2bb2ai_2 _15616_ (.A1_N(_06493_),
    .A2_N(_06496_),
    .B1(_06431_),
    .B2(_06432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_2 _15617_ (.A(_06497_),
    .B(_06498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06499_));
 sky130_fd_sc_hd__a21o_2 _15618_ (.A1(_06455_),
    .A2(_06459_),
    .B1(_06499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06500_));
 sky130_fd_sc_hd__nand3_2 _15619_ (.A(_06455_),
    .B(_06459_),
    .C(_06499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_2 _15620_ (.A(_06500_),
    .B(_06501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06502_));
 sky130_fd_sc_hd__a2bb2o_2 _15621_ (.A1_N(_06426_),
    .A2_N(_06456_),
    .B1(_06500_),
    .B2(_06501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06503_));
 sky130_fd_sc_hd__nand3_2 _15622_ (.A(_06500_),
    .B(_06501_),
    .C(_06458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06504_));
 sky130_fd_sc_hd__o311a_2 _15623_ (.A1(_06426_),
    .A2(_06456_),
    .A3(_06502_),
    .B1(_06503_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00343_));
 sky130_fd_sc_hd__nand2_2 _15624_ (.A(\a_l[0] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06505_));
 sky130_fd_sc_hd__a31o_2 _15625_ (.A1(\a_l[0] ),
    .A2(_06466_),
    .A3(\b_h[5] ),
    .B1(_06468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06506_));
 sky130_fd_sc_hd__a21o_2 _15626_ (.A1(\a_l[0] ),
    .A2(\b_h[6] ),
    .B1(_06506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06507_));
 sky130_fd_sc_hd__and3_2 _15627_ (.A(_06506_),
    .B(\b_h[6] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06508_));
 sky130_fd_sc_hd__nand3_2 _15628_ (.A(_06506_),
    .B(\b_h[6] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06509_));
 sky130_fd_sc_hd__nand2_2 _15629_ (.A(_06507_),
    .B(_06509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06510_));
 sky130_fd_sc_hd__inv_2 _15630_ (.A(_06510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_2 _15631_ (.A(_06472_),
    .B(_06490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06512_));
 sky130_fd_sc_hd__a32oi_2 _15632_ (.A1(_06474_),
    .A2(_06483_),
    .A3(_06484_),
    .B1(_06490_),
    .B2(_06472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06513_));
 sky130_fd_sc_hd__a32o_2 _15633_ (.A1(_06474_),
    .A2(_06483_),
    .A3(_06484_),
    .B1(_06490_),
    .B2(_06472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06514_));
 sky130_fd_sc_hd__o21ai_2 _15634_ (.A1(_06475_),
    .A2(_06478_),
    .B1(_06481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06515_));
 sky130_fd_sc_hd__nand2_2 _15635_ (.A(_06479_),
    .B(_06486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06516_));
 sky130_fd_sc_hd__nor2_2 _15636_ (.A(_09210_),
    .B(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06517_));
 sky130_fd_sc_hd__nand2_2 _15637_ (.A(\a_l[5] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06518_));
 sky130_fd_sc_hd__nand2_2 _15638_ (.A(\a_l[3] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06519_));
 sky130_fd_sc_hd__nand2_2 _15639_ (.A(\a_l[4] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06520_));
 sky130_fd_sc_hd__nand2_2 _15640_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06521_));
 sky130_fd_sc_hd__nand4_2 _15641_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06522_));
 sky130_fd_sc_hd__a22oi_2 _15642_ (.A1(\a_l[4] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06523_));
 sky130_fd_sc_hd__nand2_2 _15643_ (.A(_06519_),
    .B(_06520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06524_));
 sky130_fd_sc_hd__o21ai_2 _15644_ (.A1(_06440_),
    .A2(_06521_),
    .B1(_06524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_2 _15645_ (.A(_06525_),
    .B(_06517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06526_));
 sky130_fd_sc_hd__o21ai_2 _15646_ (.A1(_06440_),
    .A2(_06521_),
    .B1(_06518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06527_));
 sky130_fd_sc_hd__o211ai_2 _15647_ (.A1(_06527_),
    .A2(_06523_),
    .B1(_06516_),
    .C1(_06526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06528_));
 sky130_fd_sc_hd__a41o_2 _15648_ (.A1(\a_l[3] ),
    .A2(\a_l[4] ),
    .A3(\b_h[2] ),
    .A4(\b_h[3] ),
    .B1(_06518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06529_));
 sky130_fd_sc_hd__o311a_2 _15649_ (.A1(_09188_),
    .A2(_09199_),
    .A3(_06440_),
    .B1(_06517_),
    .C1(_06524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06530_));
 sky130_fd_sc_hd__o2bb2ai_2 _15650_ (.A1_N(_06522_),
    .A2_N(_06524_),
    .B1(_09210_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_2 _15651_ (.A(_06531_),
    .B(_06515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06532_));
 sky130_fd_sc_hd__o211ai_2 _15652_ (.A1(_06523_),
    .A2(_06529_),
    .B1(_06515_),
    .C1(_06531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06533_));
 sky130_fd_sc_hd__and2_2 _15653_ (.A(\a_l[1] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06534_));
 sky130_fd_sc_hd__nand2_2 _15654_ (.A(\a_l[1] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06535_));
 sky130_fd_sc_hd__nand2_2 _15655_ (.A(\a_l[2] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_2 _15656_ (.A(\a_l[6] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06537_));
 sky130_fd_sc_hd__o21a_2 _15657_ (.A1(_09231_),
    .A2(_09526_),
    .B1(_06536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06538_));
 sky130_fd_sc_hd__nand2_2 _15658_ (.A(_06536_),
    .B(_06537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06539_));
 sky130_fd_sc_hd__nand4_2 _15659_ (.A(\a_l[2] ),
    .B(\a_l[6] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06540_));
 sky130_fd_sc_hd__a21oi_2 _15660_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06541_));
 sky130_fd_sc_hd__a21o_2 _15661_ (.A1(_06539_),
    .A2(_06540_),
    .B1(_06534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_2 _15662_ (.A1(_06536_),
    .A2(_06537_),
    .B1(_06535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06543_));
 sky130_fd_sc_hd__o21ai_2 _15663_ (.A1(_06536_),
    .A2(_06537_),
    .B1(_06543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06544_));
 sky130_fd_sc_hd__a21oi_2 _15664_ (.A1(_06540_),
    .A2(_06543_),
    .B1(_06541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_2 _15665_ (.A(_06542_),
    .B(_06544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06546_));
 sky130_fd_sc_hd__o2111ai_2 _15666_ (.A1(_06530_),
    .A2(_06532_),
    .B1(_06542_),
    .C1(_06544_),
    .D1(_06528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06547_));
 sky130_fd_sc_hd__a21o_2 _15667_ (.A1(_06528_),
    .A2(_06533_),
    .B1(_06545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06548_));
 sky130_fd_sc_hd__a21oi_2 _15668_ (.A1(_06528_),
    .A2(_06533_),
    .B1(_06546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06549_));
 sky130_fd_sc_hd__a21o_2 _15669_ (.A1(_06528_),
    .A2(_06533_),
    .B1(_06546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06550_));
 sky130_fd_sc_hd__nand3_2 _15670_ (.A(_06528_),
    .B(_06533_),
    .C(_06546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06551_));
 sky130_fd_sc_hd__o211ai_2 _15671_ (.A1(_06482_),
    .A2(_06488_),
    .B1(_06512_),
    .C1(_06551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06552_));
 sky130_fd_sc_hd__nand3_2 _15672_ (.A(_06550_),
    .B(_06551_),
    .C(_06513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06553_));
 sky130_fd_sc_hd__a21oi_2 _15673_ (.A1(_06550_),
    .A2(_06551_),
    .B1(_06513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06554_));
 sky130_fd_sc_hd__nand3_2 _15674_ (.A(_06514_),
    .B(_06547_),
    .C(_06548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06555_));
 sky130_fd_sc_hd__o21bai_2 _15675_ (.A1(_06549_),
    .A2(_06552_),
    .B1_N(_06510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06556_));
 sky130_fd_sc_hd__a22o_2 _15676_ (.A1(_06507_),
    .A2(_06509_),
    .B1(_06553_),
    .B2(_06555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06557_));
 sky130_fd_sc_hd__o211ai_2 _15677_ (.A1(_06552_),
    .A2(_06549_),
    .B1(_06510_),
    .C1(_06555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06558_));
 sky130_fd_sc_hd__a21o_2 _15678_ (.A1(_06553_),
    .A2(_06555_),
    .B1(_06510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06559_));
 sky130_fd_sc_hd__o21ai_2 _15679_ (.A1(_06554_),
    .A2(_06556_),
    .B1(_06557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_2 _15680_ (.A(_06493_),
    .B(_06433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_2 _15681_ (.A(_06496_),
    .B(_06561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06562_));
 sky130_fd_sc_hd__inv_2 _15682_ (.A(_06562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06563_));
 sky130_fd_sc_hd__o211a_2 _15683_ (.A1(_06554_),
    .A2(_06556_),
    .B1(_06562_),
    .C1(_06557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06564_));
 sky130_fd_sc_hd__o211ai_2 _15684_ (.A1(_06554_),
    .A2(_06556_),
    .B1(_06562_),
    .C1(_06557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06565_));
 sky130_fd_sc_hd__nand4_2 _15685_ (.A(_06496_),
    .B(_06558_),
    .C(_06559_),
    .D(_06561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_2 _15686_ (.A(_06565_),
    .B(_06566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06567_));
 sky130_fd_sc_hd__a2bb2o_2 _15687_ (.A1_N(_06455_),
    .A2_N(_06499_),
    .B1(_06565_),
    .B2(_06566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06568_));
 sky130_fd_sc_hd__a211oi_2 _15688_ (.A1(_06560_),
    .A2(_06563_),
    .B1(_06455_),
    .C1(_06499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06569_));
 sky130_fd_sc_hd__nand4b_2 _15689_ (.A_N(_06455_),
    .B(_06497_),
    .C(_06498_),
    .D(_06566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06570_));
 sky130_fd_sc_hd__nand2_2 _15690_ (.A(_06568_),
    .B(_06570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06571_));
 sky130_fd_sc_hd__or2_2 _15691_ (.A(_06459_),
    .B(_06499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06572_));
 sky130_fd_sc_hd__a21oi_2 _15692_ (.A1(_06504_),
    .A2(_06572_),
    .B1(_06571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06573_));
 sky130_fd_sc_hd__a31o_2 _15693_ (.A1(_06504_),
    .A2(_06571_),
    .A3(_06572_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06574_));
 sky130_fd_sc_hd__nor2_2 _15694_ (.A(_06573_),
    .B(_06574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_2 _15695_ (.A(_06555_),
    .B(_06556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06575_));
 sky130_fd_sc_hd__a21oi_2 _15696_ (.A1(_06511_),
    .A2(_06553_),
    .B1(_06554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06576_));
 sky130_fd_sc_hd__nand2_2 _15697_ (.A(\a_l[1] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06577_));
 sky130_fd_sc_hd__and4_2 _15698_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06578_));
 sky130_fd_sc_hd__a22oi_2 _15699_ (.A1(\a_l[1] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06579_));
 sky130_fd_sc_hd__o31a_2 _15700_ (.A1(_09231_),
    .A2(_09526_),
    .A3(_06536_),
    .B1(_06535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06580_));
 sky130_fd_sc_hd__a2111oi_2 _15701_ (.A1(_06535_),
    .A2(_06540_),
    .B1(_06578_),
    .C1(_06579_),
    .D1(_06538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06581_));
 sky130_fd_sc_hd__or4_2 _15702_ (.A(_06538_),
    .B(_06578_),
    .C(_06579_),
    .D(_06580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06582_));
 sky130_fd_sc_hd__o22a_2 _15703_ (.A1(_06578_),
    .A2(_06579_),
    .B1(_06580_),
    .B2(_06538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06583_));
 sky130_fd_sc_hd__nor2_2 _15704_ (.A(_06581_),
    .B(_06583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06584_));
 sky130_fd_sc_hd__a21boi_2 _15705_ (.A1(_06528_),
    .A2(_06545_),
    .B1_N(_06533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06585_));
 sky130_fd_sc_hd__o2bb2ai_2 _15706_ (.A1_N(_06545_),
    .A2_N(_06528_),
    .B1(_06532_),
    .B2(_06530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06586_));
 sky130_fd_sc_hd__nand2_2 _15707_ (.A(\a_l[2] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06587_));
 sky130_fd_sc_hd__nand2_2 _15708_ (.A(\a_l[3] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2_2 _15709_ (.A(\a_l[7] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06589_));
 sky130_fd_sc_hd__a22oi_2 _15710_ (.A1(\a_l[7] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06590_));
 sky130_fd_sc_hd__nand2_2 _15711_ (.A(_06588_),
    .B(_06589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06591_));
 sky130_fd_sc_hd__nand4_2 _15712_ (.A(\a_l[3] ),
    .B(\a_l[7] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06592_));
 sky130_fd_sc_hd__a22oi_2 _15713_ (.A1(\a_l[2] ),
    .A2(\b_h[5] ),
    .B1(_06591_),
    .B2(_06592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06593_));
 sky130_fd_sc_hd__a21oi_2 _15714_ (.A1(_06588_),
    .A2(_06589_),
    .B1(_06587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06594_));
 sky130_fd_sc_hd__and4_2 _15715_ (.A(_06591_),
    .B(_06592_),
    .C(\a_l[2] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06595_));
 sky130_fd_sc_hd__a21oi_2 _15716_ (.A1(_06592_),
    .A2(_06594_),
    .B1(_06593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06596_));
 sky130_fd_sc_hd__a21o_2 _15717_ (.A1(_06518_),
    .A2(_06522_),
    .B1(_06523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06597_));
 sky130_fd_sc_hd__a21oi_2 _15718_ (.A1(_06518_),
    .A2(_06522_),
    .B1(_06523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06598_));
 sky130_fd_sc_hd__and2_2 _15719_ (.A(\a_l[6] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06599_));
 sky130_fd_sc_hd__nand2_2 _15720_ (.A(\a_l[6] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06600_));
 sky130_fd_sc_hd__nand2_2 _15721_ (.A(\a_l[4] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06601_));
 sky130_fd_sc_hd__nand2_2 _15722_ (.A(\a_l[5] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06602_));
 sky130_fd_sc_hd__a22oi_2 _15723_ (.A1(\a_l[5] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06603_));
 sky130_fd_sc_hd__nand2_2 _15724_ (.A(_06601_),
    .B(_06602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06604_));
 sky130_fd_sc_hd__nand2_2 _15725_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06605_));
 sky130_fd_sc_hd__and4_2 _15726_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06606_));
 sky130_fd_sc_hd__nand4_2 _15727_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06607_));
 sky130_fd_sc_hd__nand2_2 _15728_ (.A(_06604_),
    .B(_06607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06608_));
 sky130_fd_sc_hd__a21oi_2 _15729_ (.A1(_06604_),
    .A2(_06607_),
    .B1(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06609_));
 sky130_fd_sc_hd__a22o_2 _15730_ (.A1(\a_l[6] ),
    .A2(\b_h[1] ),
    .B1(_06604_),
    .B2(_06607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06610_));
 sky130_fd_sc_hd__o211ai_2 _15731_ (.A1(_06440_),
    .A2(_06605_),
    .B1(_06599_),
    .C1(_06604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06611_));
 sky130_fd_sc_hd__o221ai_2 _15732_ (.A1(_09231_),
    .A2(_09581_),
    .B1(_06440_),
    .B2(_06605_),
    .C1(_06604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_2 _15733_ (.A(_06608_),
    .B(_06599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06613_));
 sky130_fd_sc_hd__nand3_2 _15734_ (.A(_06613_),
    .B(_06597_),
    .C(_06612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06614_));
 sky130_fd_sc_hd__nand2_2 _15735_ (.A(_06598_),
    .B(_06611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06615_));
 sky130_fd_sc_hd__nand4_2 _15736_ (.A(_06524_),
    .B(_06527_),
    .C(_06610_),
    .D(_06611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06616_));
 sky130_fd_sc_hd__o21ai_2 _15737_ (.A1(_06609_),
    .A2(_06615_),
    .B1(_06614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06617_));
 sky130_fd_sc_hd__o21ai_2 _15738_ (.A1(_06593_),
    .A2(_06595_),
    .B1(_06617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06618_));
 sky130_fd_sc_hd__o211ai_2 _15739_ (.A1(_06609_),
    .A2(_06615_),
    .B1(_06596_),
    .C1(_06614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06619_));
 sky130_fd_sc_hd__inv_2 _15740_ (.A(_06619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06620_));
 sky130_fd_sc_hd__o211ai_2 _15741_ (.A1(_06593_),
    .A2(_06595_),
    .B1(_06614_),
    .C1(_06616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06621_));
 sky130_fd_sc_hd__nand2_2 _15742_ (.A(_06617_),
    .B(_06596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06622_));
 sky130_fd_sc_hd__and3_2 _15743_ (.A(_06622_),
    .B(_06585_),
    .C(_06621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06623_));
 sky130_fd_sc_hd__nand3_2 _15744_ (.A(_06622_),
    .B(_06585_),
    .C(_06621_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06624_));
 sky130_fd_sc_hd__nand2_2 _15745_ (.A(_06586_),
    .B(_06618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06625_));
 sky130_fd_sc_hd__nand3_2 _15746_ (.A(_06586_),
    .B(_06618_),
    .C(_06619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06626_));
 sky130_fd_sc_hd__nand2_2 _15747_ (.A(_06624_),
    .B(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06627_));
 sky130_fd_sc_hd__o21ai_2 _15748_ (.A1(_06581_),
    .A2(_06583_),
    .B1(_06627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06628_));
 sky130_fd_sc_hd__o211ai_2 _15749_ (.A1(_06620_),
    .A2(_06625_),
    .B1(_06624_),
    .C1(_06584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06629_));
 sky130_fd_sc_hd__a31oi_2 _15750_ (.A1(_06586_),
    .A2(_06618_),
    .A3(_06619_),
    .B1(_06584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06630_));
 sky130_fd_sc_hd__o21ai_2 _15751_ (.A1(_06581_),
    .A2(_06583_),
    .B1(_06626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_2 _15752_ (.A(_06630_),
    .B(_06624_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06632_));
 sky130_fd_sc_hd__nand2_2 _15753_ (.A(_06627_),
    .B(_06584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06633_));
 sky130_fd_sc_hd__o211ai_2 _15754_ (.A1(_06631_),
    .A2(_06623_),
    .B1(_06576_),
    .C1(_06633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06634_));
 sky130_fd_sc_hd__a21oi_2 _15755_ (.A1(_06632_),
    .A2(_06633_),
    .B1(_06576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06635_));
 sky130_fd_sc_hd__nand3_2 _15756_ (.A(_06628_),
    .B(_06629_),
    .C(_06575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06636_));
 sky130_fd_sc_hd__nand2_2 _15757_ (.A(_06634_),
    .B(_06636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06637_));
 sky130_fd_sc_hd__nand3_2 _15758_ (.A(_06509_),
    .B(_06634_),
    .C(_06636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06638_));
 sky130_fd_sc_hd__nand2_2 _15759_ (.A(_06637_),
    .B(_06508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06639_));
 sky130_fd_sc_hd__a21o_2 _15760_ (.A1(_06634_),
    .A2(_06636_),
    .B1(_06508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06640_));
 sky130_fd_sc_hd__nand3_2 _15761_ (.A(_06634_),
    .B(_06636_),
    .C(_06508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_2 _15762_ (.A(_06638_),
    .B(_06639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06642_));
 sky130_fd_sc_hd__o211ai_2 _15763_ (.A1(_06560_),
    .A2(_06563_),
    .B1(_06638_),
    .C1(_06639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06643_));
 sky130_fd_sc_hd__nand3_2 _15764_ (.A(_06640_),
    .B(_06641_),
    .C(_06564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06644_));
 sky130_fd_sc_hd__nand2_2 _15765_ (.A(_06643_),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06645_));
 sky130_fd_sc_hd__o21a_2 _15766_ (.A1(_06567_),
    .A2(_06572_),
    .B1(_06570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06646_));
 sky130_fd_sc_hd__nand2_2 _15767_ (.A(_06645_),
    .B(_06646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06647_));
 sky130_fd_sc_hd__mux2_1 _15768_ (.A0(_06643_),
    .A1(_06645_),
    .S(_06646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06648_));
 sky130_fd_sc_hd__nand3b_2 _15769_ (.A_N(_06504_),
    .B(_06568_),
    .C(_06570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06649_));
 sky130_fd_sc_hd__a21oi_2 _15770_ (.A1(_06645_),
    .A2(_06646_),
    .B1(_06649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06650_));
 sky130_fd_sc_hd__and4_2 _15771_ (.A(_06501_),
    .B(_06568_),
    .C(_06647_),
    .D(_06460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06651_));
 sky130_fd_sc_hd__a211oi_2 _15772_ (.A1(_06648_),
    .A2(_06649_),
    .B1(_06650_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00345_));
 sky130_fd_sc_hd__a31oi_2 _15773_ (.A1(_06576_),
    .A2(_06632_),
    .A3(_06633_),
    .B1(_06509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06652_));
 sky130_fd_sc_hd__a21o_2 _15774_ (.A1(_06508_),
    .A2(_06634_),
    .B1(_06635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06653_));
 sky130_fd_sc_hd__o2bb2ai_2 _15775_ (.A1_N(_06584_),
    .A2_N(_06624_),
    .B1(_06620_),
    .B2(_06625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06654_));
 sky130_fd_sc_hd__o21ai_2 _15776_ (.A1(_06587_),
    .A2(_06590_),
    .B1(_06592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06655_));
 sky130_fd_sc_hd__o21a_2 _15777_ (.A1(_06587_),
    .A2(_06590_),
    .B1(_06592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06656_));
 sky130_fd_sc_hd__nand2_2 _15778_ (.A(\a_l[0] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06657_));
 sky130_fd_sc_hd__nand2_2 _15779_ (.A(\a_l[2] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06658_));
 sky130_fd_sc_hd__nand2_2 _15780_ (.A(_06577_),
    .B(_06658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06659_));
 sky130_fd_sc_hd__and4_2 _15781_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06660_));
 sky130_fd_sc_hd__nand4_2 _15782_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06661_));
 sky130_fd_sc_hd__nand4_2 _15783_ (.A(_06659_),
    .B(_06661_),
    .C(\a_l[0] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06662_));
 sky130_fd_sc_hd__a22o_2 _15784_ (.A1(\a_l[0] ),
    .A2(\b_h[8] ),
    .B1(_06659_),
    .B2(_06661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06663_));
 sky130_fd_sc_hd__nand3_2 _15785_ (.A(_06663_),
    .B(_06655_),
    .C(_06662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06664_));
 sky130_fd_sc_hd__o211ai_2 _15786_ (.A1(_09166_),
    .A2(_09613_),
    .B1(_06659_),
    .C1(_06661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06665_));
 sky130_fd_sc_hd__a21o_2 _15787_ (.A1(_06659_),
    .A2(_06661_),
    .B1(_06657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06666_));
 sky130_fd_sc_hd__nand3_2 _15788_ (.A(_06656_),
    .B(_06665_),
    .C(_06666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06667_));
 sky130_fd_sc_hd__a21boi_2 _15789_ (.A1(_06664_),
    .A2(_06667_),
    .B1_N(_06578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06668_));
 sky130_fd_sc_hd__o211a_2 _15790_ (.A1(_06505_),
    .A2(_06577_),
    .B1(_06664_),
    .C1(_06667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06669_));
 sky130_fd_sc_hd__o2bb2ai_2 _15791_ (.A1_N(_06664_),
    .A2_N(_06667_),
    .B1(_06505_),
    .B2(_06577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06670_));
 sky130_fd_sc_hd__nand3_2 _15792_ (.A(_06667_),
    .B(_06578_),
    .C(_06664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06671_));
 sky130_fd_sc_hd__nand2_2 _15793_ (.A(_06670_),
    .B(_06671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06672_));
 sky130_fd_sc_hd__o2bb2ai_2 _15794_ (.A1_N(_06596_),
    .A2_N(_06614_),
    .B1(_06615_),
    .B2(_06609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06673_));
 sky130_fd_sc_hd__a2bb2oi_2 _15795_ (.A1_N(_06609_),
    .A2_N(_06615_),
    .B1(_06596_),
    .B2(_06614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06674_));
 sky130_fd_sc_hd__a21o_2 _15796_ (.A1(_06600_),
    .A2(_06607_),
    .B1(_06603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06675_));
 sky130_fd_sc_hd__a21oi_2 _15797_ (.A1(_06600_),
    .A2(_06607_),
    .B1(_06603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06676_));
 sky130_fd_sc_hd__nand2_2 _15798_ (.A(\a_l[7] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_2 _15799_ (.A(\a_l[5] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06678_));
 sky130_fd_sc_hd__nand2_2 _15800_ (.A(\a_l[6] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06679_));
 sky130_fd_sc_hd__nand2_2 _15801_ (.A(_06678_),
    .B(_06679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06680_));
 sky130_fd_sc_hd__nand2_2 _15802_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06681_));
 sky130_fd_sc_hd__and4_2 _15803_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06682_));
 sky130_fd_sc_hd__nand4_2 _15804_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06683_));
 sky130_fd_sc_hd__o2bb2a_2 _15805_ (.A1_N(_06680_),
    .A2_N(_06683_),
    .B1(_09242_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06684_));
 sky130_fd_sc_hd__o2bb2ai_2 _15806_ (.A1_N(_06680_),
    .A2_N(_06683_),
    .B1(_09242_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06685_));
 sky130_fd_sc_hd__o2111ai_2 _15807_ (.A1(_06440_),
    .A2(_06681_),
    .B1(\a_l[7] ),
    .C1(\b_h[1] ),
    .D1(_06680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06686_));
 sky130_fd_sc_hd__o221ai_2 _15808_ (.A1(_09242_),
    .A2(_09581_),
    .B1(_06440_),
    .B2(_06681_),
    .C1(_06680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06687_));
 sky130_fd_sc_hd__a21o_2 _15809_ (.A1(_06680_),
    .A2(_06683_),
    .B1(_06677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06688_));
 sky130_fd_sc_hd__nand3_2 _15810_ (.A(_06688_),
    .B(_06675_),
    .C(_06687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06689_));
 sky130_fd_sc_hd__o211ai_2 _15811_ (.A1(_06599_),
    .A2(_06606_),
    .B1(_06686_),
    .C1(_06604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06690_));
 sky130_fd_sc_hd__nand3_2 _15812_ (.A(_06676_),
    .B(_06685_),
    .C(_06686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06691_));
 sky130_fd_sc_hd__nand2_2 _15813_ (.A(\a_l[3] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_2 _15814_ (.A(\a_l[4] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06693_));
 sky130_fd_sc_hd__nand2_2 _15815_ (.A(\a_l[8] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06694_));
 sky130_fd_sc_hd__a22oi_2 _15816_ (.A1(\a_l[8] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_2 _15817_ (.A(_06693_),
    .B(_06694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06696_));
 sky130_fd_sc_hd__nand4_2 _15818_ (.A(\a_l[4] ),
    .B(\a_l[8] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06697_));
 sky130_fd_sc_hd__o2bb2a_2 _15819_ (.A1_N(_06696_),
    .A2_N(_06697_),
    .B1(_09188_),
    .B2(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06698_));
 sky130_fd_sc_hd__and4_2 _15820_ (.A(_06696_),
    .B(_06697_),
    .C(\a_l[3] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06699_));
 sky130_fd_sc_hd__a21oi_2 _15821_ (.A1(_06696_),
    .A2(_06697_),
    .B1(_06692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06700_));
 sky130_fd_sc_hd__a21o_2 _15822_ (.A1(_06696_),
    .A2(_06697_),
    .B1(_06692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06701_));
 sky130_fd_sc_hd__and3_2 _15823_ (.A(_06692_),
    .B(_06696_),
    .C(_06697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06702_));
 sky130_fd_sc_hd__o211ai_2 _15824_ (.A1(_09188_),
    .A2(_09602_),
    .B1(_06696_),
    .C1(_06697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06703_));
 sky130_fd_sc_hd__nand2_2 _15825_ (.A(_06701_),
    .B(_06703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06704_));
 sky130_fd_sc_hd__nand4_2 _15826_ (.A(_06689_),
    .B(_06691_),
    .C(_06701_),
    .D(_06703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06705_));
 sky130_fd_sc_hd__o2bb2ai_2 _15827_ (.A1_N(_06689_),
    .A2_N(_06691_),
    .B1(_06700_),
    .B2(_06702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06706_));
 sky130_fd_sc_hd__o2bb2ai_2 _15828_ (.A1_N(_06689_),
    .A2_N(_06691_),
    .B1(_06698_),
    .B2(_06699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06707_));
 sky130_fd_sc_hd__o211ai_2 _15829_ (.A1(_06700_),
    .A2(_06702_),
    .B1(_06689_),
    .C1(_06691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06708_));
 sky130_fd_sc_hd__nand3_2 _15830_ (.A(_06674_),
    .B(_06705_),
    .C(_06706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06709_));
 sky130_fd_sc_hd__nand3_2 _15831_ (.A(_06707_),
    .B(_06708_),
    .C(_06673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06710_));
 sky130_fd_sc_hd__nand2_2 _15832_ (.A(_06709_),
    .B(_06710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_2 _15833_ (.A(_06710_),
    .B(_06672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06712_));
 sky130_fd_sc_hd__and3_2 _15834_ (.A(_06709_),
    .B(_06710_),
    .C(_06672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06713_));
 sky130_fd_sc_hd__nand3_2 _15835_ (.A(_06709_),
    .B(_06710_),
    .C(_06672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06714_));
 sky130_fd_sc_hd__o21ai_2 _15836_ (.A1(_06668_),
    .A2(_06669_),
    .B1(_06711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06715_));
 sky130_fd_sc_hd__o211ai_2 _15837_ (.A1(_06668_),
    .A2(_06669_),
    .B1(_06709_),
    .C1(_06710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06716_));
 sky130_fd_sc_hd__nand2_2 _15838_ (.A(_06711_),
    .B(_06672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06717_));
 sky130_fd_sc_hd__o21ai_2 _15839_ (.A1(_06623_),
    .A2(_06630_),
    .B1(_06715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06718_));
 sky130_fd_sc_hd__a2bb2oi_2 _15840_ (.A1_N(_06623_),
    .A2_N(_06630_),
    .B1(_06716_),
    .B2(_06717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06719_));
 sky130_fd_sc_hd__o211ai_2 _15841_ (.A1(_06623_),
    .A2(_06630_),
    .B1(_06714_),
    .C1(_06715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06720_));
 sky130_fd_sc_hd__nand3_2 _15842_ (.A(_06717_),
    .B(_06654_),
    .C(_06716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06721_));
 sky130_fd_sc_hd__a21o_2 _15843_ (.A1(_06720_),
    .A2(_06721_),
    .B1(_06581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06722_));
 sky130_fd_sc_hd__o211ai_2 _15844_ (.A1(_06713_),
    .A2(_06718_),
    .B1(_06721_),
    .C1(_06581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06723_));
 sky130_fd_sc_hd__o211ai_2 _15845_ (.A1(_06713_),
    .A2(_06718_),
    .B1(_06721_),
    .C1(_06582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06724_));
 sky130_fd_sc_hd__a21o_2 _15846_ (.A1(_06720_),
    .A2(_06721_),
    .B1(_06582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06725_));
 sky130_fd_sc_hd__a21oi_2 _15847_ (.A1(_06722_),
    .A2(_06723_),
    .B1(_06653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06726_));
 sky130_fd_sc_hd__nand4_2 _15848_ (.A(_06636_),
    .B(_06641_),
    .C(_06724_),
    .D(_06725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06727_));
 sky130_fd_sc_hd__a2bb2oi_2 _15849_ (.A1_N(_06635_),
    .A2_N(_06652_),
    .B1(_06724_),
    .B2(_06725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06728_));
 sky130_fd_sc_hd__o211ai_2 _15850_ (.A1(_06635_),
    .A2(_06652_),
    .B1(_06722_),
    .C1(_06723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_2 _15851_ (.A(_06727_),
    .B(_06729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06730_));
 sky130_fd_sc_hd__nand2_2 _15852_ (.A(_06643_),
    .B(_06569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06731_));
 sky130_fd_sc_hd__nand2_2 _15853_ (.A(_06570_),
    .B(_06644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06732_));
 sky130_fd_sc_hd__a21o_2 _15854_ (.A1(_06644_),
    .A2(_06731_),
    .B1(_06730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06733_));
 sky130_fd_sc_hd__o211ai_2 _15855_ (.A1(_06642_),
    .A2(_06564_),
    .B1(_06732_),
    .C1(_06730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06734_));
 sky130_fd_sc_hd__nand4_2 _15856_ (.A(_06644_),
    .B(_06727_),
    .C(_06729_),
    .D(_06731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_2 _15857_ (.A(_06734_),
    .B(_06735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06736_));
 sky130_fd_sc_hd__and4b_2 _15858_ (.A_N(_06572_),
    .B(_06642_),
    .C(_06565_),
    .D(_06566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06737_));
 sky130_fd_sc_hd__o2bb2ai_2 _15859_ (.A1_N(_06734_),
    .A2_N(_06735_),
    .B1(_06737_),
    .B2(_06650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06738_));
 sky130_fd_sc_hd__o21ai_2 _15860_ (.A1(_06651_),
    .A2(_06737_),
    .B1(_06736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06739_));
 sky130_fd_sc_hd__o311a_2 _15861_ (.A1(_06651_),
    .A2(_06736_),
    .A3(_06737_),
    .B1(_06738_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00346_));
 sky130_fd_sc_hd__o41a_2 _15862_ (.A1(_06538_),
    .A2(_06578_),
    .A3(_06579_),
    .A4(_06580_),
    .B1(_06721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06740_));
 sky130_fd_sc_hd__o2bb2ai_2 _15863_ (.A1_N(_06582_),
    .A2_N(_06721_),
    .B1(_06713_),
    .B2(_06718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06741_));
 sky130_fd_sc_hd__a21oi_2 _15864_ (.A1(_06582_),
    .A2(_06721_),
    .B1(_06719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_2 _15865_ (.A(\a_l[0] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06743_));
 sky130_fd_sc_hd__a32oi_2 _15866_ (.A1(_06655_),
    .A2(_06662_),
    .A3(_06663_),
    .B1(_06667_),
    .B2(_06578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06744_));
 sky130_fd_sc_hd__nor2_2 _15867_ (.A(_06743_),
    .B(_06744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06745_));
 sky130_fd_sc_hd__or3_2 _15868_ (.A(_09166_),
    .B(_09624_),
    .C(_06744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06746_));
 sky130_fd_sc_hd__o21a_2 _15869_ (.A1(_09166_),
    .A2(_09624_),
    .B1(_06744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06747_));
 sky130_fd_sc_hd__nor2_2 _15870_ (.A(_06745_),
    .B(_06747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06748_));
 sky130_fd_sc_hd__nand2_2 _15871_ (.A(_06709_),
    .B(_06712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06749_));
 sky130_fd_sc_hd__o2bb2ai_2 _15872_ (.A1_N(_06704_),
    .A2_N(_06689_),
    .B1(_06684_),
    .B2(_06690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06750_));
 sky130_fd_sc_hd__a21boi_2 _15873_ (.A1(_06689_),
    .A2(_06704_),
    .B1_N(_06691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06751_));
 sky130_fd_sc_hd__a21oi_2 _15874_ (.A1(_06678_),
    .A2(_06679_),
    .B1(_06677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06752_));
 sky130_fd_sc_hd__nand2_2 _15875_ (.A(_06677_),
    .B(_06683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06753_));
 sky130_fd_sc_hd__nand2_2 _15876_ (.A(_06680_),
    .B(_06753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06754_));
 sky130_fd_sc_hd__a31o_2 _15877_ (.A1(\a_l[7] ),
    .A2(_06680_),
    .A3(\b_h[1] ),
    .B1(_06682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06755_));
 sky130_fd_sc_hd__nand2_2 _15878_ (.A(\a_l[8] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06756_));
 sky130_fd_sc_hd__nand2_2 _15879_ (.A(\a_l[6] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_2 _15880_ (.A(\a_l[7] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06758_));
 sky130_fd_sc_hd__a22oi_2 _15881_ (.A1(\a_l[7] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_2 _15882_ (.A(_06757_),
    .B(_06758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_2 _15883_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06761_));
 sky130_fd_sc_hd__nand4_2 _15884_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06762_));
 sky130_fd_sc_hd__nand4_2 _15885_ (.A(_06760_),
    .B(_06762_),
    .C(\a_l[8] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06763_));
 sky130_fd_sc_hd__o2bb2ai_2 _15886_ (.A1_N(_06760_),
    .A2_N(_06762_),
    .B1(_09253_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06764_));
 sky130_fd_sc_hd__o211ai_2 _15887_ (.A1(_09253_),
    .A2(_09581_),
    .B1(_06760_),
    .C1(_06762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06765_));
 sky130_fd_sc_hd__a21o_2 _15888_ (.A1(_06760_),
    .A2(_06762_),
    .B1(_06756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06766_));
 sky130_fd_sc_hd__nand2_2 _15889_ (.A(_06765_),
    .B(_06766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06767_));
 sky130_fd_sc_hd__o211a_2 _15890_ (.A1(_06682_),
    .A2(_06752_),
    .B1(_06763_),
    .C1(_06764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06768_));
 sky130_fd_sc_hd__o211ai_2 _15891_ (.A1(_06682_),
    .A2(_06752_),
    .B1(_06763_),
    .C1(_06764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06769_));
 sky130_fd_sc_hd__nand3_2 _15892_ (.A(_06766_),
    .B(_06754_),
    .C(_06765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06770_));
 sky130_fd_sc_hd__nand2_2 _15893_ (.A(\a_l[4] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06771_));
 sky130_fd_sc_hd__nand2_2 _15894_ (.A(\a_l[9] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06772_));
 sky130_fd_sc_hd__a22oi_2 _15895_ (.A1(\a_l[9] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06773_));
 sky130_fd_sc_hd__nand2_2 _15896_ (.A(_06467_),
    .B(_06772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06774_));
 sky130_fd_sc_hd__nand4_2 _15897_ (.A(\a_l[5] ),
    .B(\a_l[9] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06775_));
 sky130_fd_sc_hd__a22oi_2 _15898_ (.A1(\a_l[4] ),
    .A2(\b_h[5] ),
    .B1(_06774_),
    .B2(_06775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06776_));
 sky130_fd_sc_hd__and4_2 _15899_ (.A(_06774_),
    .B(_06775_),
    .C(\a_l[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06777_));
 sky130_fd_sc_hd__and3_2 _15900_ (.A(_06771_),
    .B(_06774_),
    .C(_06775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06778_));
 sky130_fd_sc_hd__o211ai_2 _15901_ (.A1(_09199_),
    .A2(_09602_),
    .B1(_06774_),
    .C1(_06775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06779_));
 sky130_fd_sc_hd__a21oi_2 _15902_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06780_));
 sky130_fd_sc_hd__a21o_2 _15903_ (.A1(_06774_),
    .A2(_06775_),
    .B1(_06771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06781_));
 sky130_fd_sc_hd__o211ai_2 _15904_ (.A1(_06776_),
    .A2(_06777_),
    .B1(_06769_),
    .C1(_06770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06782_));
 sky130_fd_sc_hd__o2bb2ai_2 _15905_ (.A1_N(_06769_),
    .A2_N(_06770_),
    .B1(_06778_),
    .B2(_06780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06783_));
 sky130_fd_sc_hd__nand3_2 _15906_ (.A(_06751_),
    .B(_06782_),
    .C(_06783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06784_));
 sky130_fd_sc_hd__o211ai_2 _15907_ (.A1(_06778_),
    .A2(_06780_),
    .B1(_06769_),
    .C1(_06770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06785_));
 sky130_fd_sc_hd__o2bb2ai_2 _15908_ (.A1_N(_06769_),
    .A2_N(_06770_),
    .B1(_06776_),
    .B2(_06777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06786_));
 sky130_fd_sc_hd__nand3_2 _15909_ (.A(_06786_),
    .B(_06750_),
    .C(_06785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06787_));
 sky130_fd_sc_hd__and3_2 _15910_ (.A(_06659_),
    .B(\b_h[8] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06788_));
 sky130_fd_sc_hd__a31o_2 _15911_ (.A1(\a_l[0] ),
    .A2(_06659_),
    .A3(\b_h[8] ),
    .B1(_06660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06789_));
 sky130_fd_sc_hd__nor2_2 _15912_ (.A(_06660_),
    .B(_06788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06790_));
 sky130_fd_sc_hd__and2_2 _15913_ (.A(\a_l[1] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06791_));
 sky130_fd_sc_hd__nand2_2 _15914_ (.A(\a_l[1] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_2 _15915_ (.A(\a_l[2] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06793_));
 sky130_fd_sc_hd__nand2_2 _15916_ (.A(\a_l[3] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06794_));
 sky130_fd_sc_hd__a22oi_2 _15917_ (.A1(\a_l[3] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06795_));
 sky130_fd_sc_hd__a22o_2 _15918_ (.A1(\a_l[3] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06796_));
 sky130_fd_sc_hd__nand2_2 _15919_ (.A(\a_l[3] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06797_));
 sky130_fd_sc_hd__o2bb2ai_2 _15920_ (.A1_N(_06793_),
    .A2_N(_06794_),
    .B1(_06797_),
    .B2(_06658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06798_));
 sky130_fd_sc_hd__nand2_2 _15921_ (.A(_06792_),
    .B(_06798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06799_));
 sky130_fd_sc_hd__o211ai_2 _15922_ (.A1(_06658_),
    .A2(_06797_),
    .B1(_06791_),
    .C1(_06796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06800_));
 sky130_fd_sc_hd__o211ai_2 _15923_ (.A1(_06658_),
    .A2(_06797_),
    .B1(_06796_),
    .C1(_06792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_2 _15924_ (.A(_06798_),
    .B(_06791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06802_));
 sky130_fd_sc_hd__nand2_2 _15925_ (.A(_06692_),
    .B(_06697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06803_));
 sky130_fd_sc_hd__o21ai_2 _15926_ (.A1(_06692_),
    .A2(_06695_),
    .B1(_06697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2_2 _15927_ (.A(_06696_),
    .B(_06803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06805_));
 sky130_fd_sc_hd__nand3_2 _15928_ (.A(_06801_),
    .B(_06802_),
    .C(_06805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06806_));
 sky130_fd_sc_hd__nand3_2 _15929_ (.A(_06799_),
    .B(_06800_),
    .C(_06804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06807_));
 sky130_fd_sc_hd__a21oi_2 _15930_ (.A1(_06806_),
    .A2(_06807_),
    .B1(_06789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06808_));
 sky130_fd_sc_hd__o211a_2 _15931_ (.A1(_06660_),
    .A2(_06788_),
    .B1(_06806_),
    .C1(_06807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06809_));
 sky130_fd_sc_hd__nor2_2 _15932_ (.A(_06789_),
    .B(_06806_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_2 _15933_ (.A(_06790_),
    .B(_06807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06811_));
 sky130_fd_sc_hd__nand2_2 _15934_ (.A(_06806_),
    .B(_06811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06812_));
 sky130_fd_sc_hd__a21oi_2 _15935_ (.A1(_06806_),
    .A2(_06811_),
    .B1(_06810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06813_));
 sky130_fd_sc_hd__and4_2 _15936_ (.A(_06789_),
    .B(_06799_),
    .C(_06800_),
    .D(_06804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06814_));
 sky130_fd_sc_hd__nor2_2 _15937_ (.A(_06808_),
    .B(_06809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06815_));
 sky130_fd_sc_hd__a21oi_2 _15938_ (.A1(_06784_),
    .A2(_06787_),
    .B1(_06815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06816_));
 sky130_fd_sc_hd__nand2_2 _15939_ (.A(_06784_),
    .B(_06815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06817_));
 sky130_fd_sc_hd__nand3_2 _15940_ (.A(_06784_),
    .B(_06815_),
    .C(_06787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06818_));
 sky130_fd_sc_hd__o2bb2ai_2 _15941_ (.A1_N(_06784_),
    .A2_N(_06787_),
    .B1(_06813_),
    .B2(_06814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06819_));
 sky130_fd_sc_hd__o211ai_2 _15942_ (.A1(_06808_),
    .A2(_06809_),
    .B1(_06784_),
    .C1(_06787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06820_));
 sky130_fd_sc_hd__nand3_2 _15943_ (.A(_06709_),
    .B(_06712_),
    .C(_06818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06821_));
 sky130_fd_sc_hd__a21oi_2 _15944_ (.A1(_06819_),
    .A2(_06820_),
    .B1(_06749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06822_));
 sky130_fd_sc_hd__nand3_2 _15945_ (.A(_06749_),
    .B(_06819_),
    .C(_06820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06823_));
 sky130_fd_sc_hd__o21ai_2 _15946_ (.A1(_06816_),
    .A2(_06821_),
    .B1(_06823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_2 _15947_ (.A(_06823_),
    .B(_06748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06825_));
 sky130_fd_sc_hd__o211a_2 _15948_ (.A1(_06816_),
    .A2(_06821_),
    .B1(_06823_),
    .C1(_06748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06826_));
 sky130_fd_sc_hd__o211ai_2 _15949_ (.A1(_06816_),
    .A2(_06821_),
    .B1(_06823_),
    .C1(_06748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06827_));
 sky130_fd_sc_hd__o21ai_2 _15950_ (.A1(_06745_),
    .A2(_06747_),
    .B1(_06824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06828_));
 sky130_fd_sc_hd__nand2_2 _15951_ (.A(_06824_),
    .B(_06748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06829_));
 sky130_fd_sc_hd__o221ai_2 _15952_ (.A1(_06745_),
    .A2(_06747_),
    .B1(_06816_),
    .B2(_06821_),
    .C1(_06823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06830_));
 sky130_fd_sc_hd__nand2_2 _15953_ (.A(_06742_),
    .B(_06828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06831_));
 sky130_fd_sc_hd__o211ai_2 _15954_ (.A1(_06825_),
    .A2(_06822_),
    .B1(_06742_),
    .C1(_06828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06832_));
 sky130_fd_sc_hd__inv_2 _15955_ (.A(_06832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06833_));
 sky130_fd_sc_hd__a2bb2oi_2 _15956_ (.A1_N(_06719_),
    .A2_N(_06740_),
    .B1(_06827_),
    .B2(_06828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06834_));
 sky130_fd_sc_hd__nand3_2 _15957_ (.A(_06829_),
    .B(_06830_),
    .C(_06741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06835_));
 sky130_fd_sc_hd__nand2_2 _15958_ (.A(_06832_),
    .B(_06835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_2 _15959_ (.A(_06729_),
    .B(_06836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06837_));
 sky130_fd_sc_hd__nor2_2 _15960_ (.A(_06644_),
    .B(_06726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06838_));
 sky130_fd_sc_hd__o211ai_2 _15961_ (.A1(_06644_),
    .A2(_06726_),
    .B1(_06729_),
    .C1(_06836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06839_));
 sky130_fd_sc_hd__nand2_2 _15962_ (.A(_06837_),
    .B(_06838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06840_));
 sky130_fd_sc_hd__and3_2 _15963_ (.A(_06728_),
    .B(_06832_),
    .C(_06835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06841_));
 sky130_fd_sc_hd__o211ai_2 _15964_ (.A1(_06729_),
    .A2(_06836_),
    .B1(_06839_),
    .C1(_06840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06842_));
 sky130_fd_sc_hd__o31a_2 _15965_ (.A1(_06570_),
    .A2(_06645_),
    .A3(_06730_),
    .B1(_06739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06843_));
 sky130_fd_sc_hd__o21a_2 _15966_ (.A1(_06842_),
    .A2(_06843_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06844_));
 sky130_fd_sc_hd__a21boi_2 _15967_ (.A1(_06842_),
    .A2(_06843_),
    .B1_N(_06844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00347_));
 sky130_fd_sc_hd__o22ai_2 _15968_ (.A1(_06733_),
    .A2(_06836_),
    .B1(_06842_),
    .B2(_06738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06845_));
 sky130_fd_sc_hd__o2bb2ai_2 _15969_ (.A1_N(_06748_),
    .A2_N(_06823_),
    .B1(_06821_),
    .B2(_06816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06846_));
 sky130_fd_sc_hd__or3_2 _15970_ (.A(_09624_),
    .B(_09635_),
    .C(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06847_));
 sky130_fd_sc_hd__o2bb2a_2 _15971_ (.A1_N(\a_l[1] ),
    .A2_N(\b_h[9] ),
    .B1(_09635_),
    .B2(_09166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06848_));
 sky130_fd_sc_hd__a31o_2 _15972_ (.A1(\b_h[9] ),
    .A2(\b_h[10] ),
    .A3(_06401_),
    .B1(_06848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06849_));
 sky130_fd_sc_hd__nor2_2 _15973_ (.A(_06812_),
    .B(_06849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06850_));
 sky130_fd_sc_hd__inv_2 _15974_ (.A(_06850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06851_));
 sky130_fd_sc_hd__and2_2 _15975_ (.A(_06812_),
    .B(_06849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06852_));
 sky130_fd_sc_hd__nor2_2 _15976_ (.A(_06850_),
    .B(_06852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06853_));
 sky130_fd_sc_hd__nand2_2 _15977_ (.A(_06787_),
    .B(_06817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06854_));
 sky130_fd_sc_hd__a21boi_2 _15978_ (.A1(_06784_),
    .A2(_06815_),
    .B1_N(_06787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06855_));
 sky130_fd_sc_hd__a32oi_2 _15979_ (.A1(_06766_),
    .A2(_06754_),
    .A3(_06765_),
    .B1(_06779_),
    .B2(_06781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06856_));
 sky130_fd_sc_hd__o21ai_2 _15980_ (.A1(_06776_),
    .A2(_06777_),
    .B1(_06769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06857_));
 sky130_fd_sc_hd__o21ai_2 _15981_ (.A1(_06755_),
    .A2(_06767_),
    .B1(_06857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06858_));
 sky130_fd_sc_hd__o21ai_2 _15982_ (.A1(_06756_),
    .A2(_06759_),
    .B1(_06762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06859_));
 sky130_fd_sc_hd__o21a_2 _15983_ (.A1(_06756_),
    .A2(_06759_),
    .B1(_06762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06860_));
 sky130_fd_sc_hd__nand2_2 _15984_ (.A(\a_l[9] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06861_));
 sky130_fd_sc_hd__nand2_2 _15985_ (.A(\a_l[7] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06862_));
 sky130_fd_sc_hd__nand2_2 _15986_ (.A(\a_l[8] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06863_));
 sky130_fd_sc_hd__a22oi_2 _15987_ (.A1(\a_l[8] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06864_));
 sky130_fd_sc_hd__nand2_2 _15988_ (.A(_06862_),
    .B(_06863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06865_));
 sky130_fd_sc_hd__nand2_2 _15989_ (.A(\a_l[8] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06866_));
 sky130_fd_sc_hd__nand2_2 _15990_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06867_));
 sky130_fd_sc_hd__nor2_2 _15991_ (.A(_06440_),
    .B(_06867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06868_));
 sky130_fd_sc_hd__nand4_2 _15992_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06869_));
 sky130_fd_sc_hd__o221ai_2 _15993_ (.A1(_09275_),
    .A2(_09581_),
    .B1(_06440_),
    .B2(_06867_),
    .C1(_06865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06870_));
 sky130_fd_sc_hd__o21bai_2 _15994_ (.A1(_06864_),
    .A2(_06868_),
    .B1_N(_06861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06871_));
 sky130_fd_sc_hd__o2111ai_2 _15995_ (.A1(_06440_),
    .A2(_06867_),
    .B1(\a_l[9] ),
    .C1(\b_h[1] ),
    .D1(_06865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06872_));
 sky130_fd_sc_hd__o21ai_2 _15996_ (.A1(_06864_),
    .A2(_06868_),
    .B1(_06861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06873_));
 sky130_fd_sc_hd__nand3_2 _15997_ (.A(_06873_),
    .B(_06859_),
    .C(_06872_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06874_));
 sky130_fd_sc_hd__nand3_2 _15998_ (.A(_06860_),
    .B(_06870_),
    .C(_06871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06875_));
 sky130_fd_sc_hd__and2_2 _15999_ (.A(\a_l[5] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06876_));
 sky130_fd_sc_hd__nand2_2 _16000_ (.A(\a_l[6] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06877_));
 sky130_fd_sc_hd__nand2_2 _16001_ (.A(\a_l[10] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06878_));
 sky130_fd_sc_hd__nand2_2 _16002_ (.A(_06877_),
    .B(_06878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06879_));
 sky130_fd_sc_hd__nand2_2 _16003_ (.A(\a_l[10] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06880_));
 sky130_fd_sc_hd__and4_2 _16004_ (.A(\a_l[6] ),
    .B(\a_l[10] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06881_));
 sky130_fd_sc_hd__nand4_2 _16005_ (.A(\a_l[6] ),
    .B(\a_l[10] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06882_));
 sky130_fd_sc_hd__a21oi_2 _16006_ (.A1(_06879_),
    .A2(_06882_),
    .B1(_06876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06883_));
 sky130_fd_sc_hd__o211a_2 _16007_ (.A1(_06537_),
    .A2(_06880_),
    .B1(_06876_),
    .C1(_06879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06884_));
 sky130_fd_sc_hd__a211oi_2 _16008_ (.A1(_06879_),
    .A2(_06882_),
    .B1(_09210_),
    .C1(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06885_));
 sky130_fd_sc_hd__o221a_2 _16009_ (.A1(_09210_),
    .A2(_09602_),
    .B1(_06537_),
    .B2(_06880_),
    .C1(_06879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06886_));
 sky130_fd_sc_hd__nor2_2 _16010_ (.A(_06883_),
    .B(_06884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06887_));
 sky130_fd_sc_hd__o2bb2ai_2 _16011_ (.A1_N(_06874_),
    .A2_N(_06875_),
    .B1(_06885_),
    .B2(_06886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06888_));
 sky130_fd_sc_hd__o211ai_2 _16012_ (.A1(_06883_),
    .A2(_06884_),
    .B1(_06874_),
    .C1(_06875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06889_));
 sky130_fd_sc_hd__inv_2 _16013_ (.A(_06889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06890_));
 sky130_fd_sc_hd__o211ai_2 _16014_ (.A1(_06885_),
    .A2(_06886_),
    .B1(_06874_),
    .C1(_06875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06891_));
 sky130_fd_sc_hd__o2bb2ai_2 _16015_ (.A1_N(_06874_),
    .A2_N(_06875_),
    .B1(_06883_),
    .B2(_06884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06892_));
 sky130_fd_sc_hd__o211a_2 _16016_ (.A1(_06768_),
    .A2(_06856_),
    .B1(_06891_),
    .C1(_06892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06893_));
 sky130_fd_sc_hd__o211ai_2 _16017_ (.A1(_06768_),
    .A2(_06856_),
    .B1(_06891_),
    .C1(_06892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06894_));
 sky130_fd_sc_hd__a21o_2 _16018_ (.A1(_06771_),
    .A2(_06775_),
    .B1(_06773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06895_));
 sky130_fd_sc_hd__a21oi_2 _16019_ (.A1(_06771_),
    .A2(_06775_),
    .B1(_06773_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06896_));
 sky130_fd_sc_hd__nand2_2 _16020_ (.A(\a_l[2] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06897_));
 sky130_fd_sc_hd__nand2_2 _16021_ (.A(\a_l[4] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06898_));
 sky130_fd_sc_hd__a22oi_2 _16022_ (.A1(\a_l[4] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06899_));
 sky130_fd_sc_hd__nand2_2 _16023_ (.A(_06797_),
    .B(_06898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_2 _16024_ (.A(\a_l[4] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06901_));
 sky130_fd_sc_hd__nand4_2 _16025_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06902_));
 sky130_fd_sc_hd__o2bb2ai_2 _16026_ (.A1_N(_06900_),
    .A2_N(_06902_),
    .B1(_09144_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06903_));
 sky130_fd_sc_hd__o2111ai_2 _16027_ (.A1(_06794_),
    .A2(_06901_),
    .B1(\a_l[2] ),
    .C1(\b_h[8] ),
    .D1(_06900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06904_));
 sky130_fd_sc_hd__o221ai_2 _16028_ (.A1(_09144_),
    .A2(_09613_),
    .B1(_06794_),
    .B2(_06901_),
    .C1(_06900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06905_));
 sky130_fd_sc_hd__a21o_2 _16029_ (.A1(_06900_),
    .A2(_06902_),
    .B1(_06897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06906_));
 sky130_fd_sc_hd__nand3_2 _16030_ (.A(_06906_),
    .B(_06895_),
    .C(_06905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06907_));
 sky130_fd_sc_hd__nand3_2 _16031_ (.A(_06896_),
    .B(_06903_),
    .C(_06904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06908_));
 sky130_fd_sc_hd__o2bb2a_2 _16032_ (.A1_N(\a_l[1] ),
    .A2_N(\b_h[8] ),
    .B1(_06658_),
    .B2(_06797_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06909_));
 sky130_fd_sc_hd__a41o_2 _16033_ (.A1(\a_l[2] ),
    .A2(\a_l[3] ),
    .A3(\b_h[6] ),
    .A4(\b_h[7] ),
    .B1(_06791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06910_));
 sky130_fd_sc_hd__o2bb2ai_2 _16034_ (.A1_N(_06907_),
    .A2_N(_06908_),
    .B1(_06909_),
    .B2(_06795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06911_));
 sky130_fd_sc_hd__nand4_2 _16035_ (.A(_06796_),
    .B(_06907_),
    .C(_06908_),
    .D(_06910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06912_));
 sky130_fd_sc_hd__nand2_2 _16036_ (.A(_06911_),
    .B(_06912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06913_));
 sky130_fd_sc_hd__inv_2 _16037_ (.A(_06913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06914_));
 sky130_fd_sc_hd__nand2_2 _16038_ (.A(_06858_),
    .B(_06888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06915_));
 sky130_fd_sc_hd__nand3_2 _16039_ (.A(_06858_),
    .B(_06888_),
    .C(_06889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06916_));
 sky130_fd_sc_hd__inv_2 _16040_ (.A(_06916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06917_));
 sky130_fd_sc_hd__a31oi_2 _16041_ (.A1(_06858_),
    .A2(_06888_),
    .A3(_06889_),
    .B1(_06913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06918_));
 sky130_fd_sc_hd__nand4_2 _16042_ (.A(_06894_),
    .B(_06911_),
    .C(_06912_),
    .D(_06916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06919_));
 sky130_fd_sc_hd__nand2_2 _16043_ (.A(_06894_),
    .B(_06916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06920_));
 sky130_fd_sc_hd__a22o_2 _16044_ (.A1(_06911_),
    .A2(_06912_),
    .B1(_06916_),
    .B2(_06894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06921_));
 sky130_fd_sc_hd__nand2_2 _16045_ (.A(_06920_),
    .B(_06914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06922_));
 sky130_fd_sc_hd__nand2_2 _16046_ (.A(_06894_),
    .B(_06913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06923_));
 sky130_fd_sc_hd__o211ai_2 _16047_ (.A1(_06890_),
    .A2(_06915_),
    .B1(_06913_),
    .C1(_06894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06924_));
 sky130_fd_sc_hd__a22oi_2 _16048_ (.A1(_06787_),
    .A2(_06817_),
    .B1(_06922_),
    .B2(_06924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06925_));
 sky130_fd_sc_hd__nand3_2 _16049_ (.A(_06921_),
    .B(_06854_),
    .C(_06919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06926_));
 sky130_fd_sc_hd__o211ai_2 _16050_ (.A1(_06923_),
    .A2(_06917_),
    .B1(_06855_),
    .C1(_06922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06927_));
 sky130_fd_sc_hd__nand2_2 _16051_ (.A(_06926_),
    .B(_06927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06928_));
 sky130_fd_sc_hd__a21boi_2 _16052_ (.A1(_06926_),
    .A2(_06927_),
    .B1_N(_06853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06929_));
 sky130_fd_sc_hd__nand2_2 _16053_ (.A(_06928_),
    .B(_06853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06930_));
 sky130_fd_sc_hd__nand3b_2 _16054_ (.A_N(_06853_),
    .B(_06926_),
    .C(_06927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06931_));
 sky130_fd_sc_hd__nand2_2 _16055_ (.A(_06927_),
    .B(_06853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06932_));
 sky130_fd_sc_hd__a21o_2 _16056_ (.A1(_06926_),
    .A2(_06927_),
    .B1(_06853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06933_));
 sky130_fd_sc_hd__o211ai_2 _16057_ (.A1(_06925_),
    .A2(_06932_),
    .B1(_06846_),
    .C1(_06933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06934_));
 sky130_fd_sc_hd__nor3b_2 _16058_ (.A(_06846_),
    .B(_06929_),
    .C_N(_06931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06935_));
 sky130_fd_sc_hd__nand3b_2 _16059_ (.A_N(_06846_),
    .B(_06930_),
    .C(_06931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06936_));
 sky130_fd_sc_hd__a21o_2 _16060_ (.A1(_06934_),
    .A2(_06936_),
    .B1(_06746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06937_));
 sky130_fd_sc_hd__o211ai_2 _16061_ (.A1(_06743_),
    .A2(_06744_),
    .B1(_06934_),
    .C1(_06936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06938_));
 sky130_fd_sc_hd__and3_2 _16062_ (.A(_06936_),
    .B(_06745_),
    .C(_06934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06939_));
 sky130_fd_sc_hd__o2bb2ai_2 _16063_ (.A1_N(_06934_),
    .A2_N(_06936_),
    .B1(_06743_),
    .B2(_06744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06940_));
 sky130_fd_sc_hd__nand2_2 _16064_ (.A(_06937_),
    .B(_06938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06941_));
 sky130_fd_sc_hd__a32oi_2 _16065_ (.A1(_06742_),
    .A2(_06827_),
    .A3(_06828_),
    .B1(_06728_),
    .B2(_06835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06942_));
 sky130_fd_sc_hd__o22ai_2 _16066_ (.A1(_06826_),
    .A2(_06831_),
    .B1(_06729_),
    .B2(_06834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2_2 _16067_ (.A(_06940_),
    .B(_06943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06944_));
 sky130_fd_sc_hd__a31o_2 _16068_ (.A1(_06745_),
    .A2(_06934_),
    .A3(_06936_),
    .B1(_06944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06945_));
 sky130_fd_sc_hd__nand3_2 _16069_ (.A(_06937_),
    .B(_06938_),
    .C(_06942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06946_));
 sky130_fd_sc_hd__a21oi_2 _16070_ (.A1(_06945_),
    .A2(_06946_),
    .B1(_06845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06947_));
 sky130_fd_sc_hd__and3_2 _16071_ (.A(_06845_),
    .B(_06945_),
    .C(_06946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06948_));
 sky130_fd_sc_hd__nor3_2 _16072_ (.A(rst),
    .B(_06947_),
    .C(_06948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00348_));
 sky130_fd_sc_hd__a21oi_2 _16073_ (.A1(_06937_),
    .A2(_06938_),
    .B1(_06832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06949_));
 sky130_fd_sc_hd__a21oi_2 _16074_ (.A1(_06746_),
    .A2(_06934_),
    .B1(_06935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06950_));
 sky130_fd_sc_hd__a21oi_2 _16075_ (.A1(_06927_),
    .A2(_06853_),
    .B1(_06925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06951_));
 sky130_fd_sc_hd__nand2_2 _16076_ (.A(_06926_),
    .B(_06932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06952_));
 sky130_fd_sc_hd__o2bb2ai_2 _16077_ (.A1_N(_06894_),
    .A2_N(_06913_),
    .B1(_06915_),
    .B2(_06890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06953_));
 sky130_fd_sc_hd__a31o_2 _16078_ (.A1(_06911_),
    .A2(_06912_),
    .A3(_06916_),
    .B1(_06893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06954_));
 sky130_fd_sc_hd__o21ai_2 _16079_ (.A1(_06876_),
    .A2(_06881_),
    .B1(_06879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06955_));
 sky130_fd_sc_hd__a31o_2 _16080_ (.A1(\a_l[5] ),
    .A2(_06879_),
    .A3(\b_h[5] ),
    .B1(_06881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06956_));
 sky130_fd_sc_hd__nand2_2 _16081_ (.A(\a_l[3] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06957_));
 sky130_fd_sc_hd__nand2_2 _16082_ (.A(\a_l[5] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06958_));
 sky130_fd_sc_hd__a22oi_2 _16083_ (.A1(\a_l[5] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06959_));
 sky130_fd_sc_hd__nand2_2 _16084_ (.A(_06901_),
    .B(_06958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06960_));
 sky130_fd_sc_hd__nand2_2 _16085_ (.A(\a_l[5] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06961_));
 sky130_fd_sc_hd__nand4_2 _16086_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06962_));
 sky130_fd_sc_hd__a22o_2 _16087_ (.A1(\a_l[3] ),
    .A2(\b_h[8] ),
    .B1(_06960_),
    .B2(_06962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06963_));
 sky130_fd_sc_hd__o2111ai_2 _16088_ (.A1(_06898_),
    .A2(_06961_),
    .B1(\a_l[3] ),
    .C1(\b_h[8] ),
    .D1(_06960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06964_));
 sky130_fd_sc_hd__o221ai_2 _16089_ (.A1(_09188_),
    .A2(_09613_),
    .B1(_06898_),
    .B2(_06961_),
    .C1(_06960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06965_));
 sky130_fd_sc_hd__a21o_2 _16090_ (.A1(_06960_),
    .A2(_06962_),
    .B1(_06957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06966_));
 sky130_fd_sc_hd__and3_2 _16091_ (.A(_06966_),
    .B(_06955_),
    .C(_06965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06967_));
 sky130_fd_sc_hd__nand3_2 _16092_ (.A(_06955_),
    .B(_06965_),
    .C(_06966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06968_));
 sky130_fd_sc_hd__nand3_2 _16093_ (.A(_06956_),
    .B(_06963_),
    .C(_06964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06969_));
 sky130_fd_sc_hd__o22a_2 _16094_ (.A1(_09144_),
    .A2(_09613_),
    .B1(_06794_),
    .B2(_06901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06970_));
 sky130_fd_sc_hd__a21oi_2 _16095_ (.A1(_06897_),
    .A2(_06902_),
    .B1(_06899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06971_));
 sky130_fd_sc_hd__o2bb2ai_2 _16096_ (.A1_N(_06968_),
    .A2_N(_06969_),
    .B1(_06970_),
    .B2(_06899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06972_));
 sky130_fd_sc_hd__nand3_2 _16097_ (.A(_06968_),
    .B(_06969_),
    .C(_06971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06973_));
 sky130_fd_sc_hd__nand2_2 _16098_ (.A(_06972_),
    .B(_06973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_2 _16099_ (.A(_06875_),
    .B(_06887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06975_));
 sky130_fd_sc_hd__a21boi_2 _16100_ (.A1(_06875_),
    .A2(_06887_),
    .B1_N(_06874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06976_));
 sky130_fd_sc_hd__nand2_2 _16101_ (.A(_06874_),
    .B(_06975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06977_));
 sky130_fd_sc_hd__o21ai_2 _16102_ (.A1(_06861_),
    .A2(_06864_),
    .B1(_06869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06978_));
 sky130_fd_sc_hd__o22a_2 _16103_ (.A1(_06440_),
    .A2(_06867_),
    .B1(_06861_),
    .B2(_06864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06979_));
 sky130_fd_sc_hd__nand2_2 _16104_ (.A(\a_l[10] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06980_));
 sky130_fd_sc_hd__nand2_2 _16105_ (.A(\a_l[9] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06981_));
 sky130_fd_sc_hd__a22oi_2 _16106_ (.A1(\a_l[9] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06982_));
 sky130_fd_sc_hd__nand2_2 _16107_ (.A(_06866_),
    .B(_06981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06983_));
 sky130_fd_sc_hd__nor2_2 _16108_ (.A(_09253_),
    .B(_09275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06984_));
 sky130_fd_sc_hd__nand2_2 _16109_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06985_));
 sky130_fd_sc_hd__nand4_2 _16110_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06986_));
 sky130_fd_sc_hd__a21o_2 _16111_ (.A1(_06983_),
    .A2(_06986_),
    .B1(_06980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06987_));
 sky130_fd_sc_hd__o211ai_2 _16112_ (.A1(_09286_),
    .A2(_09581_),
    .B1(_06983_),
    .C1(_06986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06988_));
 sky130_fd_sc_hd__and3_2 _16113_ (.A(_06979_),
    .B(_06987_),
    .C(_06988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06989_));
 sky130_fd_sc_hd__nand3_2 _16114_ (.A(_06979_),
    .B(_06987_),
    .C(_06988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06990_));
 sky130_fd_sc_hd__nand4_2 _16115_ (.A(_06983_),
    .B(_06986_),
    .C(\a_l[10] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06991_));
 sky130_fd_sc_hd__o2bb2ai_2 _16116_ (.A1_N(_06983_),
    .A2_N(_06986_),
    .B1(_09286_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06992_));
 sky130_fd_sc_hd__and3_2 _16117_ (.A(_06992_),
    .B(_06978_),
    .C(_06991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06993_));
 sky130_fd_sc_hd__nand3_2 _16118_ (.A(_06992_),
    .B(_06978_),
    .C(_06991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06994_));
 sky130_fd_sc_hd__nand2_2 _16119_ (.A(\a_l[6] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06995_));
 sky130_fd_sc_hd__nand2_2 _16120_ (.A(\a_l[7] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06996_));
 sky130_fd_sc_hd__nand2_2 _16121_ (.A(\a_l[11] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06997_));
 sky130_fd_sc_hd__a22o_2 _16122_ (.A1(\a_l[11] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_06998_));
 sky130_fd_sc_hd__nand2_2 _16123_ (.A(\a_l[11] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_06999_));
 sky130_fd_sc_hd__and4_2 _16124_ (.A(\a_l[7] ),
    .B(\a_l[11] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07000_));
 sky130_fd_sc_hd__nand4_2 _16125_ (.A(\a_l[7] ),
    .B(\a_l[11] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07001_));
 sky130_fd_sc_hd__a22oi_2 _16126_ (.A1(\a_l[6] ),
    .A2(\b_h[5] ),
    .B1(_06998_),
    .B2(_07001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07002_));
 sky130_fd_sc_hd__and4_2 _16127_ (.A(_06998_),
    .B(_07001_),
    .C(\a_l[6] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07003_));
 sky130_fd_sc_hd__o21ai_2 _16128_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_06995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07004_));
 sky130_fd_sc_hd__o221a_2 _16129_ (.A1(_09231_),
    .A2(_09602_),
    .B1(_06589_),
    .B2(_06999_),
    .C1(_06998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07005_));
 sky130_fd_sc_hd__a21o_2 _16130_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_07004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07006_));
 sky130_fd_sc_hd__a21oi_2 _16131_ (.A1(_06998_),
    .A2(_07001_),
    .B1(_06995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07007_));
 sky130_fd_sc_hd__a21o_2 _16132_ (.A1(_06998_),
    .A2(_07001_),
    .B1(_06995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07008_));
 sky130_fd_sc_hd__nand4_2 _16133_ (.A(_06990_),
    .B(_06994_),
    .C(_07006_),
    .D(_07008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07009_));
 sky130_fd_sc_hd__o2bb2ai_2 _16134_ (.A1_N(_06990_),
    .A2_N(_06994_),
    .B1(_07005_),
    .B2(_07007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07010_));
 sky130_fd_sc_hd__o2bb2ai_2 _16135_ (.A1_N(_06990_),
    .A2_N(_06994_),
    .B1(_07002_),
    .B2(_07003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07011_));
 sky130_fd_sc_hd__a32oi_2 _16136_ (.A1(_06979_),
    .A2(_06987_),
    .A3(_06988_),
    .B1(_07006_),
    .B2(_07008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07012_));
 sky130_fd_sc_hd__o211ai_2 _16137_ (.A1(_07005_),
    .A2(_07007_),
    .B1(_06990_),
    .C1(_06994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07013_));
 sky130_fd_sc_hd__nand3_2 _16138_ (.A(_06977_),
    .B(_07011_),
    .C(_07013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07014_));
 sky130_fd_sc_hd__a21oi_2 _16139_ (.A1(_07011_),
    .A2(_07013_),
    .B1(_06977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07015_));
 sky130_fd_sc_hd__nand3_2 _16140_ (.A(_07010_),
    .B(_06976_),
    .C(_07009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07016_));
 sky130_fd_sc_hd__nand2_2 _16141_ (.A(_07014_),
    .B(_07016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07017_));
 sky130_fd_sc_hd__nand4_2 _16142_ (.A(_06972_),
    .B(_06973_),
    .C(_07014_),
    .D(_07016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07018_));
 sky130_fd_sc_hd__nand2_2 _16143_ (.A(_07017_),
    .B(_06974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07019_));
 sky130_fd_sc_hd__a21o_2 _16144_ (.A1(_07014_),
    .A2(_07016_),
    .B1(_06974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07020_));
 sky130_fd_sc_hd__nand3_2 _16145_ (.A(_06974_),
    .B(_07014_),
    .C(_07016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07021_));
 sky130_fd_sc_hd__o211ai_2 _16146_ (.A1(_06893_),
    .A2(_06918_),
    .B1(_07018_),
    .C1(_07019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07022_));
 sky130_fd_sc_hd__nand3_2 _16147_ (.A(_07020_),
    .B(_07021_),
    .C(_06953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07023_));
 sky130_fd_sc_hd__inv_2 _16148_ (.A(_07023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07024_));
 sky130_fd_sc_hd__nand2_2 _16149_ (.A(_07022_),
    .B(_07023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07025_));
 sky130_fd_sc_hd__nand2_2 _16150_ (.A(\a_l[0] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07026_));
 sky130_fd_sc_hd__a22oi_2 _16151_ (.A1(\a_l[2] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07027_));
 sky130_fd_sc_hd__and4_2 _16152_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07028_));
 sky130_fd_sc_hd__o22a_2 _16153_ (.A1(_09166_),
    .A2(_09646_),
    .B1(_07027_),
    .B2(_07028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07029_));
 sky130_fd_sc_hd__nor4_2 _16154_ (.A(_09166_),
    .B(_09646_),
    .C(_07027_),
    .D(_07028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07030_));
 sky130_fd_sc_hd__o32a_2 _16155_ (.A1(_09624_),
    .A2(_09635_),
    .A3(_06402_),
    .B1(_07029_),
    .B2(_07030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07031_));
 sky130_fd_sc_hd__nor3_2 _16156_ (.A(_06847_),
    .B(_07029_),
    .C(_07030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07032_));
 sky130_fd_sc_hd__or2_2 _16157_ (.A(_07031_),
    .B(_07032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07033_));
 sky130_fd_sc_hd__and2_2 _16158_ (.A(_06908_),
    .B(_06912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07034_));
 sky130_fd_sc_hd__a211oi_2 _16159_ (.A1(_06908_),
    .A2(_06912_),
    .B1(_07031_),
    .C1(_07032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07035_));
 sky130_fd_sc_hd__o211a_2 _16160_ (.A1(_07031_),
    .A2(_07032_),
    .B1(_06908_),
    .C1(_06912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07036_));
 sky130_fd_sc_hd__nor2_2 _16161_ (.A(_07035_),
    .B(_07036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07037_));
 sky130_fd_sc_hd__nand2_2 _16162_ (.A(_07025_),
    .B(_07037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07038_));
 sky130_fd_sc_hd__a31oi_2 _16163_ (.A1(_06954_),
    .A2(_07018_),
    .A3(_07019_),
    .B1(_07037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07039_));
 sky130_fd_sc_hd__o211ai_2 _16164_ (.A1(_07035_),
    .A2(_07036_),
    .B1(_07022_),
    .C1(_07023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07040_));
 sky130_fd_sc_hd__o2bb2ai_2 _16165_ (.A1_N(_07022_),
    .A2_N(_07023_),
    .B1(_07035_),
    .B2(_07036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07041_));
 sky130_fd_sc_hd__nand3_2 _16166_ (.A(_07022_),
    .B(_07023_),
    .C(_07037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07042_));
 sky130_fd_sc_hd__a21oi_2 _16167_ (.A1(_07041_),
    .A2(_07042_),
    .B1(_06952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07043_));
 sky130_fd_sc_hd__nand3_2 _16168_ (.A(_07038_),
    .B(_07040_),
    .C(_06951_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07044_));
 sky130_fd_sc_hd__and3_2 _16169_ (.A(_06952_),
    .B(_07041_),
    .C(_07042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07045_));
 sky130_fd_sc_hd__nand3_2 _16170_ (.A(_06952_),
    .B(_07041_),
    .C(_07042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07046_));
 sky130_fd_sc_hd__nand3_2 _16171_ (.A(_07046_),
    .B(_06850_),
    .C(_07044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07047_));
 sky130_fd_sc_hd__inv_2 _16172_ (.A(_07047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07048_));
 sky130_fd_sc_hd__o2bb2ai_2 _16173_ (.A1_N(_07044_),
    .A2_N(_07046_),
    .B1(_06812_),
    .B2(_06849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07049_));
 sky130_fd_sc_hd__nand2_2 _16174_ (.A(_06950_),
    .B(_07049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07050_));
 sky130_fd_sc_hd__nand3_2 _16175_ (.A(_06950_),
    .B(_07047_),
    .C(_07049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07051_));
 sky130_fd_sc_hd__a21o_2 _16176_ (.A1(_07047_),
    .A2(_07049_),
    .B1(_06950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07052_));
 sky130_fd_sc_hd__a21oi_2 _16177_ (.A1(_07051_),
    .A2(_07052_),
    .B1(_06949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07053_));
 sky130_fd_sc_hd__a31o_2 _16178_ (.A1(_06833_),
    .A2(_06941_),
    .A3(_07052_),
    .B1(_07053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07054_));
 sky130_fd_sc_hd__a21oi_2 _16179_ (.A1(_06841_),
    .A2(_06941_),
    .B1(_06948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07055_));
 sky130_fd_sc_hd__a21oi_2 _16180_ (.A1(_07055_),
    .A2(_07054_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07056_));
 sky130_fd_sc_hd__o21a_2 _16181_ (.A1(_07054_),
    .A2(_07055_),
    .B1(_07056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00349_));
 sky130_fd_sc_hd__a22oi_2 _16182_ (.A1(_06841_),
    .A2(_06941_),
    .B1(_06949_),
    .B2(_07052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07057_));
 sky130_fd_sc_hd__o2111a_2 _16183_ (.A1(_06939_),
    .A2(_06944_),
    .B1(_06946_),
    .C1(_07051_),
    .D1(_07052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07058_));
 sky130_fd_sc_hd__o2bb2a_2 _16184_ (.A1_N(_07058_),
    .A2_N(_06845_),
    .B1(_07053_),
    .B2(_07057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07059_));
 sky130_fd_sc_hd__o2bb2ai_2 _16185_ (.A1_N(_07058_),
    .A2_N(_06845_),
    .B1(_07053_),
    .B2(_07057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_2 _16186_ (.A(_07023_),
    .B(_07037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07061_));
 sky130_fd_sc_hd__nand2_2 _16187_ (.A(_07022_),
    .B(_07061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07062_));
 sky130_fd_sc_hd__a31oi_2 _16188_ (.A1(_06956_),
    .A2(_06963_),
    .A3(_06964_),
    .B1(_06971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07063_));
 sky130_fd_sc_hd__nor2_2 _16189_ (.A(_06967_),
    .B(_07063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07064_));
 sky130_fd_sc_hd__o22ai_2 _16190_ (.A1(_02338_),
    .A2(_06441_),
    .B1(_07026_),
    .B2(_07027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07065_));
 sky130_fd_sc_hd__nand2_2 _16191_ (.A(\a_l[1] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07066_));
 sky130_fd_sc_hd__a22oi_2 _16192_ (.A1(\a_l[3] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07067_));
 sky130_fd_sc_hd__a22o_2 _16193_ (.A1(\a_l[3] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07068_));
 sky130_fd_sc_hd__nor2_2 _16194_ (.A(_02338_),
    .B(_06480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07069_));
 sky130_fd_sc_hd__o21ai_2 _16195_ (.A1(_07067_),
    .A2(_07069_),
    .B1(_07066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07070_));
 sky130_fd_sc_hd__a41o_2 _16196_ (.A1(\a_l[2] ),
    .A2(\a_l[3] ),
    .A3(\b_h[9] ),
    .A4(\b_h[10] ),
    .B1(_07066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07071_));
 sky130_fd_sc_hd__o211ai_2 _16197_ (.A1(_07067_),
    .A2(_07069_),
    .B1(\a_l[1] ),
    .C1(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07072_));
 sky130_fd_sc_hd__o211ai_2 _16198_ (.A1(_02338_),
    .A2(_06480_),
    .B1(_07066_),
    .C1(_07068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07073_));
 sky130_fd_sc_hd__nand3b_2 _16199_ (.A_N(_07065_),
    .B(_07072_),
    .C(_07073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07074_));
 sky130_fd_sc_hd__o211a_2 _16200_ (.A1(_07071_),
    .A2(_07067_),
    .B1(_07065_),
    .C1(_07070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07075_));
 sky130_fd_sc_hd__o211ai_2 _16201_ (.A1(_07071_),
    .A2(_07067_),
    .B1(_07065_),
    .C1(_07070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07076_));
 sky130_fd_sc_hd__nor2_2 _16202_ (.A(_09166_),
    .B(_09657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07077_));
 sky130_fd_sc_hd__nand2_2 _16203_ (.A(\a_l[0] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07078_));
 sky130_fd_sc_hd__nand4_2 _16204_ (.A(_07074_),
    .B(_07076_),
    .C(\a_l[0] ),
    .D(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07079_));
 sky130_fd_sc_hd__a22o_2 _16205_ (.A1(\a_l[0] ),
    .A2(\b_h[12] ),
    .B1(_07074_),
    .B2(_07076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07080_));
 sky130_fd_sc_hd__nand3_2 _16206_ (.A(_07080_),
    .B(_07064_),
    .C(_07079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07081_));
 sky130_fd_sc_hd__o211ai_2 _16207_ (.A1(_09166_),
    .A2(_09657_),
    .B1(_07074_),
    .C1(_07076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07082_));
 sky130_fd_sc_hd__a21o_2 _16208_ (.A1(_07074_),
    .A2(_07076_),
    .B1(_07078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07083_));
 sky130_fd_sc_hd__o211ai_2 _16209_ (.A1(_06967_),
    .A2(_07063_),
    .B1(_07082_),
    .C1(_07083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07084_));
 sky130_fd_sc_hd__or4b_2 _16210_ (.A(_06847_),
    .B(_07029_),
    .C(_07030_),
    .D_N(_07084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07085_));
 sky130_fd_sc_hd__a21bo_2 _16211_ (.A1(_07081_),
    .A2(_07084_),
    .B1_N(_07032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07086_));
 sky130_fd_sc_hd__o311ai_2 _16212_ (.A1(_06847_),
    .A2(_07029_),
    .A3(_07030_),
    .B1(_07081_),
    .C1(_07084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07087_));
 sky130_fd_sc_hd__nand2_2 _16213_ (.A(_07086_),
    .B(_07087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07088_));
 sky130_fd_sc_hd__a21o_2 _16214_ (.A1(_06974_),
    .A2(_07014_),
    .B1(_07015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07089_));
 sky130_fd_sc_hd__a21oi_2 _16215_ (.A1(_06974_),
    .A2(_07014_),
    .B1(_07015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07090_));
 sky130_fd_sc_hd__o21a_2 _16216_ (.A1(_07002_),
    .A2(_07003_),
    .B1(_06994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07091_));
 sky130_fd_sc_hd__o22a_2 _16217_ (.A1(_09286_),
    .A2(_09581_),
    .B1(_06866_),
    .B2(_06981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07092_));
 sky130_fd_sc_hd__a21oi_2 _16218_ (.A1(_06980_),
    .A2(_06986_),
    .B1(_06982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07093_));
 sky130_fd_sc_hd__and2_2 _16219_ (.A(\a_l[11] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07094_));
 sky130_fd_sc_hd__nand2_2 _16220_ (.A(\a_l[11] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_2 _16221_ (.A(\a_l[9] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07096_));
 sky130_fd_sc_hd__nand2_2 _16222_ (.A(\a_l[10] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07097_));
 sky130_fd_sc_hd__a22oi_2 _16223_ (.A1(\a_l[10] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_2 _16224_ (.A(_07096_),
    .B(_07097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07099_));
 sky130_fd_sc_hd__nand2_2 _16225_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07100_));
 sky130_fd_sc_hd__nand3_2 _16226_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07101_));
 sky130_fd_sc_hd__nand4_2 _16227_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07102_));
 sky130_fd_sc_hd__a22oi_2 _16228_ (.A1(\a_l[11] ),
    .A2(\b_h[1] ),
    .B1(_07099_),
    .B2(_07102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07103_));
 sky130_fd_sc_hd__o2bb2ai_2 _16229_ (.A1_N(_07099_),
    .A2_N(_07102_),
    .B1(_09297_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07104_));
 sky130_fd_sc_hd__o211a_2 _16230_ (.A1(_09592_),
    .A2(_07101_),
    .B1(_07094_),
    .C1(_07099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07105_));
 sky130_fd_sc_hd__o2111ai_2 _16231_ (.A1(_09592_),
    .A2(_07101_),
    .B1(\b_h[1] ),
    .C1(_07099_),
    .D1(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07106_));
 sky130_fd_sc_hd__o22a_2 _16232_ (.A1(_06982_),
    .A2(_07092_),
    .B1(_07103_),
    .B2(_07105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07107_));
 sky130_fd_sc_hd__o22ai_2 _16233_ (.A1(_06982_),
    .A2(_07092_),
    .B1(_07103_),
    .B2(_07105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07108_));
 sky130_fd_sc_hd__nand3_2 _16234_ (.A(_07093_),
    .B(_07104_),
    .C(_07106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07109_));
 sky130_fd_sc_hd__nand2_2 _16235_ (.A(\a_l[7] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07110_));
 sky130_fd_sc_hd__a22oi_2 _16236_ (.A1(\a_l[12] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07111_));
 sky130_fd_sc_hd__a22o_2 _16237_ (.A1(\a_l[12] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07112_));
 sky130_fd_sc_hd__nand2_2 _16238_ (.A(\a_l[12] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07113_));
 sky130_fd_sc_hd__nand4_2 _16239_ (.A(\a_l[8] ),
    .B(\a_l[12] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07114_));
 sky130_fd_sc_hd__a22oi_2 _16240_ (.A1(\a_l[7] ),
    .A2(\b_h[5] ),
    .B1(_07112_),
    .B2(_07114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07115_));
 sky130_fd_sc_hd__a22o_2 _16241_ (.A1(\a_l[7] ),
    .A2(\b_h[5] ),
    .B1(_07112_),
    .B2(_07114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07116_));
 sky130_fd_sc_hd__and3_2 _16242_ (.A(_07114_),
    .B(\b_h[5] ),
    .C(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07117_));
 sky130_fd_sc_hd__a41o_2 _16243_ (.A1(\a_l[8] ),
    .A2(\a_l[12] ),
    .A3(\b_h[0] ),
    .A4(\b_h[4] ),
    .B1(_07110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07118_));
 sky130_fd_sc_hd__a21oi_2 _16244_ (.A1(_07112_),
    .A2(_07117_),
    .B1(_07115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07119_));
 sky130_fd_sc_hd__o21ai_2 _16245_ (.A1(_07111_),
    .A2(_07118_),
    .B1(_07116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07120_));
 sky130_fd_sc_hd__nand3_2 _16246_ (.A(_07108_),
    .B(_07119_),
    .C(_07109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07121_));
 sky130_fd_sc_hd__a21o_2 _16247_ (.A1(_07108_),
    .A2(_07109_),
    .B1(_07119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07122_));
 sky130_fd_sc_hd__and3_2 _16248_ (.A(_07108_),
    .B(_07109_),
    .C(_07120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07123_));
 sky130_fd_sc_hd__nand3_2 _16249_ (.A(_07108_),
    .B(_07109_),
    .C(_07120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07124_));
 sky130_fd_sc_hd__a21o_2 _16250_ (.A1(_07108_),
    .A2(_07109_),
    .B1(_07120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07125_));
 sky130_fd_sc_hd__o21ai_2 _16251_ (.A1(_06989_),
    .A2(_07091_),
    .B1(_07125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07126_));
 sky130_fd_sc_hd__o211ai_2 _16252_ (.A1(_06989_),
    .A2(_07091_),
    .B1(_07124_),
    .C1(_07125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07127_));
 sky130_fd_sc_hd__o211ai_2 _16253_ (.A1(_06993_),
    .A2(_07012_),
    .B1(_07121_),
    .C1(_07122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07128_));
 sky130_fd_sc_hd__nand2_2 _16254_ (.A(\a_l[6] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07129_));
 sky130_fd_sc_hd__a22o_2 _16255_ (.A1(\a_l[6] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07130_));
 sky130_fd_sc_hd__nand2_2 _16256_ (.A(\a_l[6] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07131_));
 sky130_fd_sc_hd__nand4_2 _16257_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07132_));
 sky130_fd_sc_hd__nand4_2 _16258_ (.A(_07130_),
    .B(_07132_),
    .C(\a_l[4] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07133_));
 sky130_fd_sc_hd__nand3_2 _16259_ (.A(_07129_),
    .B(\b_h[7] ),
    .C(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07134_));
 sky130_fd_sc_hd__nand3_2 _16260_ (.A(_06961_),
    .B(\b_h[6] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07135_));
 sky130_fd_sc_hd__o211ai_2 _16261_ (.A1(_09199_),
    .A2(_09613_),
    .B1(_07134_),
    .C1(_07135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07136_));
 sky130_fd_sc_hd__a21oi_2 _16262_ (.A1(_06996_),
    .A2(_06997_),
    .B1(_06995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07137_));
 sky130_fd_sc_hd__o211a_2 _16263_ (.A1(_07000_),
    .A2(_07137_),
    .B1(_07136_),
    .C1(_07133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07138_));
 sky130_fd_sc_hd__a22oi_2 _16264_ (.A1(_06998_),
    .A2(_07004_),
    .B1(_07133_),
    .B2(_07136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07139_));
 sky130_fd_sc_hd__a211o_2 _16265_ (.A1(_06901_),
    .A2(_06958_),
    .B1(_09188_),
    .C1(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07140_));
 sky130_fd_sc_hd__o32a_2 _16266_ (.A1(_09188_),
    .A2(_09613_),
    .A3(_06959_),
    .B1(_06961_),
    .B2(_06898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07141_));
 sky130_fd_sc_hd__a21oi_2 _16267_ (.A1(_06957_),
    .A2(_06962_),
    .B1(_06959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07142_));
 sky130_fd_sc_hd__o21a_2 _16268_ (.A1(_07138_),
    .A2(_07139_),
    .B1(_07142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07143_));
 sky130_fd_sc_hd__nor3_2 _16269_ (.A(_07142_),
    .B(_07139_),
    .C(_07138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07144_));
 sky130_fd_sc_hd__o21ai_2 _16270_ (.A1(_07138_),
    .A2(_07139_),
    .B1(_07141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07145_));
 sky130_fd_sc_hd__inv_2 _16271_ (.A(_07145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07146_));
 sky130_fd_sc_hd__a21o_2 _16272_ (.A1(_06962_),
    .A2(_07140_),
    .B1(_07139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07147_));
 sky130_fd_sc_hd__nor2_2 _16273_ (.A(_07138_),
    .B(_07147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07148_));
 sky130_fd_sc_hd__o21ai_2 _16274_ (.A1(_07138_),
    .A2(_07147_),
    .B1(_07145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07149_));
 sky130_fd_sc_hd__o2111ai_2 _16275_ (.A1(_07138_),
    .A2(_07147_),
    .B1(_07145_),
    .C1(_07127_),
    .D1(_07128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07150_));
 sky130_fd_sc_hd__o2bb2ai_2 _16276_ (.A1_N(_07127_),
    .A2_N(_07128_),
    .B1(_07146_),
    .B2(_07148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07151_));
 sky130_fd_sc_hd__o2bb2ai_2 _16277_ (.A1_N(_07127_),
    .A2_N(_07128_),
    .B1(_07143_),
    .B2(_07144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07152_));
 sky130_fd_sc_hd__o211ai_2 _16278_ (.A1(_07123_),
    .A2(_07126_),
    .B1(_07128_),
    .C1(_07149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07153_));
 sky130_fd_sc_hd__a21oi_2 _16279_ (.A1(_07152_),
    .A2(_07153_),
    .B1(_07089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07154_));
 sky130_fd_sc_hd__nand3_2 _16280_ (.A(_07090_),
    .B(_07150_),
    .C(_07151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07155_));
 sky130_fd_sc_hd__nand3_2 _16281_ (.A(_07089_),
    .B(_07152_),
    .C(_07153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_2 _16282_ (.A(_07155_),
    .B(_07156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07157_));
 sky130_fd_sc_hd__nand4_2 _16283_ (.A(_07086_),
    .B(_07087_),
    .C(_07155_),
    .D(_07156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07158_));
 sky130_fd_sc_hd__nand2_2 _16284_ (.A(_07157_),
    .B(_07088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07159_));
 sky130_fd_sc_hd__a32oi_2 _16285_ (.A1(_07089_),
    .A2(_07152_),
    .A3(_07153_),
    .B1(_07087_),
    .B2(_07086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07160_));
 sky130_fd_sc_hd__and3_2 _16286_ (.A(_07088_),
    .B(_07155_),
    .C(_07156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07161_));
 sky130_fd_sc_hd__nand3_2 _16287_ (.A(_07088_),
    .B(_07155_),
    .C(_07156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07162_));
 sky130_fd_sc_hd__a21o_2 _16288_ (.A1(_07155_),
    .A2(_07156_),
    .B1(_07088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07163_));
 sky130_fd_sc_hd__nand2_2 _16289_ (.A(_07163_),
    .B(_07062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07164_));
 sky130_fd_sc_hd__nand3_2 _16290_ (.A(_07163_),
    .B(_07062_),
    .C(_07162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07165_));
 sky130_fd_sc_hd__o211ai_2 _16291_ (.A1(_07024_),
    .A2(_07039_),
    .B1(_07158_),
    .C1(_07159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07166_));
 sky130_fd_sc_hd__a21oi_2 _16292_ (.A1(_07165_),
    .A2(_07166_),
    .B1(_07035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07167_));
 sky130_fd_sc_hd__o2bb2ai_2 _16293_ (.A1_N(_07165_),
    .A2_N(_07166_),
    .B1(_07033_),
    .B2(_07034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07168_));
 sky130_fd_sc_hd__and3_2 _16294_ (.A(_07165_),
    .B(_07166_),
    .C(_07035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07169_));
 sky130_fd_sc_hd__nand3_2 _16295_ (.A(_07166_),
    .B(_07035_),
    .C(_07165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07170_));
 sky130_fd_sc_hd__nor2_2 _16296_ (.A(_07167_),
    .B(_07169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2_2 _16297_ (.A(_07168_),
    .B(_07170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07172_));
 sky130_fd_sc_hd__a31oi_2 _16298_ (.A1(_06951_),
    .A2(_07038_),
    .A3(_07040_),
    .B1(_06851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07173_));
 sky130_fd_sc_hd__o21ai_2 _16299_ (.A1(_06851_),
    .A2(_07043_),
    .B1(_07046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07174_));
 sky130_fd_sc_hd__inv_2 _16300_ (.A(_07174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07175_));
 sky130_fd_sc_hd__o211a_2 _16301_ (.A1(_07045_),
    .A2(_07173_),
    .B1(_07170_),
    .C1(_07168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07176_));
 sky130_fd_sc_hd__o211ai_2 _16302_ (.A1(_07045_),
    .A2(_07173_),
    .B1(_07170_),
    .C1(_07168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07177_));
 sky130_fd_sc_hd__a21oi_2 _16303_ (.A1(_07168_),
    .A2(_07170_),
    .B1(_07174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07178_));
 sky130_fd_sc_hd__a21o_2 _16304_ (.A1(_07168_),
    .A2(_07170_),
    .B1(_07174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07179_));
 sky130_fd_sc_hd__and4b_2 _16305_ (.A_N(_07050_),
    .B(_07177_),
    .C(_07179_),
    .D(_07047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07180_));
 sky130_fd_sc_hd__nand3b_2 _16306_ (.A_N(_07051_),
    .B(_07177_),
    .C(_07179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07181_));
 sky130_fd_sc_hd__o22ai_2 _16307_ (.A1(_07050_),
    .A2(_07048_),
    .B1(_07178_),
    .B2(_07176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_2 _16308_ (.A(_07181_),
    .B(_07182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07183_));
 sky130_fd_sc_hd__and3_2 _16309_ (.A(_07060_),
    .B(_07181_),
    .C(_07182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07184_));
 sky130_fd_sc_hd__a31o_2 _16310_ (.A1(_07060_),
    .A2(_07181_),
    .A3(_07182_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07185_));
 sky130_fd_sc_hd__a21oi_2 _16311_ (.A1(_07059_),
    .A2(_07183_),
    .B1(_07185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00350_));
 sky130_fd_sc_hd__a21o_2 _16312_ (.A1(_07060_),
    .A2(_07182_),
    .B1(_07180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07186_));
 sky130_fd_sc_hd__a21oi_2 _16313_ (.A1(_07088_),
    .A2(_07156_),
    .B1(_07154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07187_));
 sky130_fd_sc_hd__o22ai_2 _16314_ (.A1(_02338_),
    .A2(_06480_),
    .B1(_07066_),
    .B2(_07067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07188_));
 sky130_fd_sc_hd__o22a_2 _16315_ (.A1(_02338_),
    .A2(_06480_),
    .B1(_07066_),
    .B2(_07067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07189_));
 sky130_fd_sc_hd__nand2_2 _16316_ (.A(\a_l[2] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2_2 _16317_ (.A(\a_l[3] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07191_));
 sky130_fd_sc_hd__nand2_2 _16318_ (.A(\a_l[4] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07192_));
 sky130_fd_sc_hd__a22oi_2 _16319_ (.A1(\a_l[4] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07193_));
 sky130_fd_sc_hd__nand2_2 _16320_ (.A(_07191_),
    .B(_07192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07194_));
 sky130_fd_sc_hd__and4_2 _16321_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07195_));
 sky130_fd_sc_hd__nand4_2 _16322_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07196_));
 sky130_fd_sc_hd__a21o_2 _16323_ (.A1(_07194_),
    .A2(_07196_),
    .B1(_07190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07197_));
 sky130_fd_sc_hd__o21ai_2 _16324_ (.A1(_07191_),
    .A2(_07192_),
    .B1(_07190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07198_));
 sky130_fd_sc_hd__o211ai_2 _16325_ (.A1(_07193_),
    .A2(_07198_),
    .B1(_07197_),
    .C1(_07189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07199_));
 sky130_fd_sc_hd__a22o_2 _16326_ (.A1(\a_l[2] ),
    .A2(\b_h[11] ),
    .B1(_07194_),
    .B2(_07196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07200_));
 sky130_fd_sc_hd__a41o_2 _16327_ (.A1(\a_l[3] ),
    .A2(\a_l[4] ),
    .A3(\b_h[9] ),
    .A4(\b_h[10] ),
    .B1(_07190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07201_));
 sky130_fd_sc_hd__o211ai_2 _16328_ (.A1(_07193_),
    .A2(_07201_),
    .B1(_07188_),
    .C1(_07200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07202_));
 sky130_fd_sc_hd__a22oi_2 _16329_ (.A1(\a_l[1] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07203_));
 sky130_fd_sc_hd__a21oi_2 _16330_ (.A1(_02588_),
    .A2(_06401_),
    .B1(_07203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07204_));
 sky130_fd_sc_hd__a31o_2 _16331_ (.A1(\a_l[1] ),
    .A2(\a_l[0] ),
    .A3(_02588_),
    .B1(_07203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07205_));
 sky130_fd_sc_hd__a21o_2 _16332_ (.A1(_07199_),
    .A2(_07202_),
    .B1(_07204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07206_));
 sky130_fd_sc_hd__nand3_2 _16333_ (.A(_07199_),
    .B(_07202_),
    .C(_07204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07207_));
 sky130_fd_sc_hd__a21o_2 _16334_ (.A1(_07199_),
    .A2(_07202_),
    .B1(_07205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07208_));
 sky130_fd_sc_hd__nand3_2 _16335_ (.A(_07199_),
    .B(_07202_),
    .C(_07205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07209_));
 sky130_fd_sc_hd__nor2_2 _16336_ (.A(_07142_),
    .B(_07138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07210_));
 sky130_fd_sc_hd__o21bai_2 _16337_ (.A1(_07139_),
    .A2(_07141_),
    .B1_N(_07138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07211_));
 sky130_fd_sc_hd__o211ai_2 _16338_ (.A1(_07139_),
    .A2(_07210_),
    .B1(_07209_),
    .C1(_07208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07212_));
 sky130_fd_sc_hd__and3_2 _16339_ (.A(_07206_),
    .B(_07211_),
    .C(_07207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07213_));
 sky130_fd_sc_hd__nand3_2 _16340_ (.A(_07206_),
    .B(_07207_),
    .C(_07211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07214_));
 sky130_fd_sc_hd__a31o_2 _16341_ (.A1(_07074_),
    .A2(\b_h[12] ),
    .A3(\a_l[0] ),
    .B1(_07075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07215_));
 sky130_fd_sc_hd__a21oi_2 _16342_ (.A1(_07074_),
    .A2(_07077_),
    .B1(_07075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07216_));
 sky130_fd_sc_hd__a21oi_2 _16343_ (.A1(_07212_),
    .A2(_07214_),
    .B1(_07215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07217_));
 sky130_fd_sc_hd__a21o_2 _16344_ (.A1(_07212_),
    .A2(_07214_),
    .B1(_07215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07218_));
 sky130_fd_sc_hd__a31oi_2 _16345_ (.A1(_07206_),
    .A2(_07211_),
    .A3(_07207_),
    .B1(_07216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07219_));
 sky130_fd_sc_hd__nand3_2 _16346_ (.A(_07212_),
    .B(_07214_),
    .C(_07215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07220_));
 sky130_fd_sc_hd__a21oi_2 _16347_ (.A1(_07212_),
    .A2(_07219_),
    .B1(_07217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07221_));
 sky130_fd_sc_hd__nand2_2 _16348_ (.A(_07218_),
    .B(_07220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07222_));
 sky130_fd_sc_hd__a2bb2oi_2 _16349_ (.A1_N(_07123_),
    .A2_N(_07126_),
    .B1(_07128_),
    .B2(_07149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07223_));
 sky130_fd_sc_hd__o2bb2ai_2 _16350_ (.A1_N(_07149_),
    .A2_N(_07128_),
    .B1(_07126_),
    .B2(_07123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07224_));
 sky130_fd_sc_hd__o21ai_2 _16351_ (.A1(_07120_),
    .A2(_07107_),
    .B1(_07109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07225_));
 sky130_fd_sc_hd__a21boi_2 _16352_ (.A1(_07108_),
    .A2(_07119_),
    .B1_N(_07109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07226_));
 sky130_fd_sc_hd__a21o_2 _16353_ (.A1(_07095_),
    .A2(_07102_),
    .B1(_07098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07227_));
 sky130_fd_sc_hd__a21oi_2 _16354_ (.A1(_07095_),
    .A2(_07102_),
    .B1(_07098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07228_));
 sky130_fd_sc_hd__nand2_2 _16355_ (.A(\a_l[12] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07229_));
 sky130_fd_sc_hd__nand2_2 _16356_ (.A(\a_l[10] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07230_));
 sky130_fd_sc_hd__nand2_2 _16357_ (.A(\a_l[11] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07231_));
 sky130_fd_sc_hd__a22oi_2 _16358_ (.A1(\a_l[11] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_2 _16359_ (.A(_07230_),
    .B(_07231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07233_));
 sky130_fd_sc_hd__nand2_2 _16360_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07234_));
 sky130_fd_sc_hd__nand4_2 _16361_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07235_));
 sky130_fd_sc_hd__a21o_2 _16362_ (.A1(_07233_),
    .A2(_07235_),
    .B1(_07229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07236_));
 sky130_fd_sc_hd__o221ai_2 _16363_ (.A1(_09319_),
    .A2(_09581_),
    .B1(_06440_),
    .B2(_07234_),
    .C1(_07233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07237_));
 sky130_fd_sc_hd__o2bb2ai_2 _16364_ (.A1_N(_07233_),
    .A2_N(_07235_),
    .B1(_09319_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07238_));
 sky130_fd_sc_hd__o2111ai_2 _16365_ (.A1(_06440_),
    .A2(_07234_),
    .B1(\a_l[12] ),
    .C1(\b_h[1] ),
    .D1(_07233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07239_));
 sky130_fd_sc_hd__nand3_2 _16366_ (.A(_07228_),
    .B(_07238_),
    .C(_07239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07240_));
 sky130_fd_sc_hd__nand3_2 _16367_ (.A(_07236_),
    .B(_07237_),
    .C(_07227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07241_));
 sky130_fd_sc_hd__a22oi_2 _16368_ (.A1(\a_l[13] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07242_));
 sky130_fd_sc_hd__a22o_2 _16369_ (.A1(\a_l[13] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07243_));
 sky130_fd_sc_hd__nand2_2 _16370_ (.A(\a_l[13] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07244_));
 sky130_fd_sc_hd__nand4_2 _16371_ (.A(\a_l[9] ),
    .B(\a_l[13] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07245_));
 sky130_fd_sc_hd__nand2_2 _16372_ (.A(\a_l[8] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07246_));
 sky130_fd_sc_hd__a22oi_2 _16373_ (.A1(\a_l[8] ),
    .A2(\b_h[5] ),
    .B1(_07243_),
    .B2(_07245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07247_));
 sky130_fd_sc_hd__a22o_2 _16374_ (.A1(\a_l[8] ),
    .A2(\b_h[5] ),
    .B1(_07243_),
    .B2(_07245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07248_));
 sky130_fd_sc_hd__a41o_2 _16375_ (.A1(\a_l[9] ),
    .A2(\a_l[13] ),
    .A3(\b_h[0] ),
    .A4(\b_h[4] ),
    .B1(_07246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07249_));
 sky130_fd_sc_hd__and4_2 _16376_ (.A(_07243_),
    .B(_07245_),
    .C(\a_l[8] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07250_));
 sky130_fd_sc_hd__o21ai_2 _16377_ (.A1(_07242_),
    .A2(_07249_),
    .B1(_07248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07251_));
 sky130_fd_sc_hd__o211ai_2 _16378_ (.A1(_07247_),
    .A2(_07250_),
    .B1(_07240_),
    .C1(_07241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07252_));
 sky130_fd_sc_hd__a21o_2 _16379_ (.A1(_07240_),
    .A2(_07241_),
    .B1(_07251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07253_));
 sky130_fd_sc_hd__o2bb2ai_2 _16380_ (.A1_N(_07240_),
    .A2_N(_07241_),
    .B1(_07247_),
    .B2(_07250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07254_));
 sky130_fd_sc_hd__o2111ai_2 _16381_ (.A1(_07242_),
    .A2(_07249_),
    .B1(_07248_),
    .C1(_07240_),
    .D1(_07241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07255_));
 sky130_fd_sc_hd__nand3_2 _16382_ (.A(_07225_),
    .B(_07254_),
    .C(_07255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07256_));
 sky130_fd_sc_hd__nand3_2 _16383_ (.A(_07226_),
    .B(_07252_),
    .C(_07253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07257_));
 sky130_fd_sc_hd__o21ai_2 _16384_ (.A1(_06961_),
    .A2(_07129_),
    .B1(_07133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07258_));
 sky130_fd_sc_hd__inv_2 _16385_ (.A(_07258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07259_));
 sky130_fd_sc_hd__nand2_2 _16386_ (.A(\a_l[7] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_2 _16387_ (.A(_07131_),
    .B(_07260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07261_));
 sky130_fd_sc_hd__nand2_2 _16388_ (.A(\a_l[7] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07262_));
 sky130_fd_sc_hd__nand4_2 _16389_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07263_));
 sky130_fd_sc_hd__nand3_2 _16390_ (.A(_07131_),
    .B(\b_h[6] ),
    .C(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07264_));
 sky130_fd_sc_hd__nand3_2 _16391_ (.A(_07260_),
    .B(\b_h[7] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07265_));
 sky130_fd_sc_hd__o211ai_2 _16392_ (.A1(_09210_),
    .A2(_09613_),
    .B1(_07264_),
    .C1(_07265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07266_));
 sky130_fd_sc_hd__nand4_2 _16393_ (.A(_07261_),
    .B(_07263_),
    .C(\a_l[5] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07267_));
 sky130_fd_sc_hd__o2bb2a_2 _16394_ (.A1_N(\a_l[7] ),
    .A2_N(\b_h[5] ),
    .B1(_06694_),
    .B2(_07113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07268_));
 sky130_fd_sc_hd__a21oi_2 _16395_ (.A1(_07110_),
    .A2(_07114_),
    .B1(_07111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07269_));
 sky130_fd_sc_hd__o2bb2ai_2 _16396_ (.A1_N(_07266_),
    .A2_N(_07267_),
    .B1(_07268_),
    .B2(_07111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07270_));
 sky130_fd_sc_hd__inv_2 _16397_ (.A(_07270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07271_));
 sky130_fd_sc_hd__nand3_2 _16398_ (.A(_07266_),
    .B(_07267_),
    .C(_07269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07272_));
 sky130_fd_sc_hd__and3_2 _16399_ (.A(_07258_),
    .B(_07270_),
    .C(_07272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07273_));
 sky130_fd_sc_hd__nand3_2 _16400_ (.A(_07258_),
    .B(_07270_),
    .C(_07272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07274_));
 sky130_fd_sc_hd__a21oi_2 _16401_ (.A1(_07270_),
    .A2(_07272_),
    .B1(_07258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07275_));
 sky130_fd_sc_hd__a21o_2 _16402_ (.A1(_07270_),
    .A2(_07272_),
    .B1(_07258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07276_));
 sky130_fd_sc_hd__a21oi_2 _16403_ (.A1(_07270_),
    .A2(_07272_),
    .B1(_07259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07277_));
 sky130_fd_sc_hd__and3_2 _16404_ (.A(_07259_),
    .B(_07270_),
    .C(_07272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07278_));
 sky130_fd_sc_hd__nand2_2 _16405_ (.A(_07274_),
    .B(_07276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07279_));
 sky130_fd_sc_hd__o211ai_2 _16406_ (.A1(_07277_),
    .A2(_07278_),
    .B1(_07256_),
    .C1(_07257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07280_));
 sky130_fd_sc_hd__o2bb2ai_2 _16407_ (.A1_N(_07256_),
    .A2_N(_07257_),
    .B1(_07273_),
    .B2(_07275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07281_));
 sky130_fd_sc_hd__o2bb2ai_2 _16408_ (.A1_N(_07256_),
    .A2_N(_07257_),
    .B1(_07277_),
    .B2(_07278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07282_));
 sky130_fd_sc_hd__nand3_2 _16409_ (.A(_07256_),
    .B(_07257_),
    .C(_07279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07283_));
 sky130_fd_sc_hd__a21oi_2 _16410_ (.A1(_07282_),
    .A2(_07283_),
    .B1(_07224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07284_));
 sky130_fd_sc_hd__nand3_2 _16411_ (.A(_07223_),
    .B(_07280_),
    .C(_07281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07285_));
 sky130_fd_sc_hd__nand3_2 _16412_ (.A(_07224_),
    .B(_07282_),
    .C(_07283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07286_));
 sky130_fd_sc_hd__nand2_2 _16413_ (.A(_07221_),
    .B(_07286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07287_));
 sky130_fd_sc_hd__a22o_2 _16414_ (.A1(_07218_),
    .A2(_07220_),
    .B1(_07285_),
    .B2(_07286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07288_));
 sky130_fd_sc_hd__o221ai_2 _16415_ (.A1(_07284_),
    .A2(_07287_),
    .B1(_07154_),
    .B2(_07160_),
    .C1(_07288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07289_));
 sky130_fd_sc_hd__nand3_2 _16416_ (.A(_07222_),
    .B(_07285_),
    .C(_07286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07290_));
 sky130_fd_sc_hd__a21o_2 _16417_ (.A1(_07285_),
    .A2(_07286_),
    .B1(_07222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07291_));
 sky130_fd_sc_hd__nand3_2 _16418_ (.A(_07187_),
    .B(_07290_),
    .C(_07291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07292_));
 sky130_fd_sc_hd__nand2_2 _16419_ (.A(_07289_),
    .B(_07292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07293_));
 sky130_fd_sc_hd__nand2_2 _16420_ (.A(_07081_),
    .B(_07085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07294_));
 sky130_fd_sc_hd__nand2_2 _16421_ (.A(_07293_),
    .B(_07294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07295_));
 sky130_fd_sc_hd__nand4_2 _16422_ (.A(_07081_),
    .B(_07085_),
    .C(_07289_),
    .D(_07292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07296_));
 sky130_fd_sc_hd__a21o_2 _16423_ (.A1(_07289_),
    .A2(_07292_),
    .B1(_07294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07297_));
 sky130_fd_sc_hd__nand3_2 _16424_ (.A(_07289_),
    .B(_07292_),
    .C(_07294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07298_));
 sky130_fd_sc_hd__o2bb2ai_2 _16425_ (.A1_N(_07035_),
    .A2_N(_07166_),
    .B1(_07164_),
    .B2(_07161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07299_));
 sky130_fd_sc_hd__a21boi_2 _16426_ (.A1(_07035_),
    .A2(_07166_),
    .B1_N(_07165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07300_));
 sky130_fd_sc_hd__nand3_2 _16427_ (.A(_07295_),
    .B(_07296_),
    .C(_07300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07301_));
 sky130_fd_sc_hd__and3_2 _16428_ (.A(_07297_),
    .B(_07298_),
    .C(_07299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07302_));
 sky130_fd_sc_hd__nand3_2 _16429_ (.A(_07297_),
    .B(_07298_),
    .C(_07299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07303_));
 sky130_fd_sc_hd__nand2_2 _16430_ (.A(_07301_),
    .B(_07303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07304_));
 sky130_fd_sc_hd__nand3_2 _16431_ (.A(_07171_),
    .B(_07301_),
    .C(_07174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07305_));
 sky130_fd_sc_hd__o2bb2ai_2 _16432_ (.A1_N(_07301_),
    .A2_N(_07303_),
    .B1(_07172_),
    .B2(_07175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07306_));
 sky130_fd_sc_hd__o41a_2 _16433_ (.A1(_07167_),
    .A2(_07169_),
    .A3(_07175_),
    .A4(_07304_),
    .B1(_07306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07307_));
 sky130_fd_sc_hd__a21oi_2 _16434_ (.A1(_07186_),
    .A2(_07307_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07308_));
 sky130_fd_sc_hd__o31a_2 _16435_ (.A1(_07180_),
    .A2(_07184_),
    .A3(_07307_),
    .B1(_07308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00351_));
 sky130_fd_sc_hd__nand2_2 _16436_ (.A(_07285_),
    .B(_07287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07309_));
 sky130_fd_sc_hd__a21boi_2 _16437_ (.A1(_07221_),
    .A2(_07286_),
    .B1_N(_07285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07310_));
 sky130_fd_sc_hd__o211a_2 _16438_ (.A1(_06961_),
    .A2(_07129_),
    .B1(_07133_),
    .C1(_07272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07311_));
 sky130_fd_sc_hd__a32o_2 _16439_ (.A1(_07266_),
    .A2(_07267_),
    .A3(_07269_),
    .B1(_07270_),
    .B2(_07258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07312_));
 sky130_fd_sc_hd__a22oi_2 _16440_ (.A1(\a_l[2] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07313_));
 sky130_fd_sc_hd__a22o_2 _16441_ (.A1(\a_l[2] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07314_));
 sky130_fd_sc_hd__and4_2 _16442_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07315_));
 sky130_fd_sc_hd__o2111a_2 _16443_ (.A1(_02589_),
    .A2(_06441_),
    .B1(\a_l[0] ),
    .C1(\b_h[14] ),
    .D1(_07314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07316_));
 sky130_fd_sc_hd__or4_2 _16444_ (.A(_09166_),
    .B(_09668_),
    .C(_07313_),
    .D(_07315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07317_));
 sky130_fd_sc_hd__o221a_2 _16445_ (.A1(_09166_),
    .A2(_09668_),
    .B1(_02589_),
    .B2(_06441_),
    .C1(_07314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07318_));
 sky130_fd_sc_hd__o211a_2 _16446_ (.A1(_07313_),
    .A2(_07315_),
    .B1(\a_l[0] ),
    .C1(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07319_));
 sky130_fd_sc_hd__nor2_2 _16447_ (.A(_07318_),
    .B(_07319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07320_));
 sky130_fd_sc_hd__a21oi_2 _16448_ (.A1(_07191_),
    .A2(_07192_),
    .B1(_07190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07321_));
 sky130_fd_sc_hd__nand2_2 _16449_ (.A(\a_l[4] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07322_));
 sky130_fd_sc_hd__nand2_2 _16450_ (.A(\a_l[5] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07323_));
 sky130_fd_sc_hd__nand2_2 _16451_ (.A(_07322_),
    .B(_07323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07324_));
 sky130_fd_sc_hd__nand3_2 _16452_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07325_));
 sky130_fd_sc_hd__nand4_2 _16453_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07326_));
 sky130_fd_sc_hd__and2_2 _16454_ (.A(\a_l[3] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07327_));
 sky130_fd_sc_hd__o2111ai_2 _16455_ (.A1(_09624_),
    .A2(_07325_),
    .B1(\b_h[11] ),
    .C1(\a_l[3] ),
    .D1(_07324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07328_));
 sky130_fd_sc_hd__o2bb2ai_2 _16456_ (.A1_N(_07324_),
    .A2_N(_07326_),
    .B1(_09188_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07329_));
 sky130_fd_sc_hd__o211a_2 _16457_ (.A1(_07195_),
    .A2(_07321_),
    .B1(_07328_),
    .C1(_07329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07330_));
 sky130_fd_sc_hd__o211ai_2 _16458_ (.A1(_07195_),
    .A2(_07321_),
    .B1(_07328_),
    .C1(_07329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07331_));
 sky130_fd_sc_hd__a22oi_2 _16459_ (.A1(_07194_),
    .A2(_07198_),
    .B1(_07328_),
    .B2(_07329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07332_));
 sky130_fd_sc_hd__a22o_2 _16460_ (.A1(_07194_),
    .A2(_07198_),
    .B1(_07328_),
    .B2(_07329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07333_));
 sky130_fd_sc_hd__o211ai_2 _16461_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07331_),
    .C1(_07333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07334_));
 sky130_fd_sc_hd__o21ai_2 _16462_ (.A1(_07330_),
    .A2(_07332_),
    .B1(_07320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07335_));
 sky130_fd_sc_hd__nand3_2 _16463_ (.A(_07320_),
    .B(_07331_),
    .C(_07333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07336_));
 sky130_fd_sc_hd__o22ai_2 _16464_ (.A1(_07318_),
    .A2(_07319_),
    .B1(_07330_),
    .B2(_07332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07337_));
 sky130_fd_sc_hd__o211ai_2 _16465_ (.A1(_07271_),
    .A2(_07311_),
    .B1(_07336_),
    .C1(_07337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07338_));
 sky130_fd_sc_hd__a21bo_2 _16466_ (.A1(_07199_),
    .A2(_07204_),
    .B1_N(_07202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07339_));
 sky130_fd_sc_hd__a21boi_2 _16467_ (.A1(_07199_),
    .A2(_07204_),
    .B1_N(_07202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07340_));
 sky130_fd_sc_hd__nand3_2 _16468_ (.A(_07335_),
    .B(_07312_),
    .C(_07334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07341_));
 sky130_fd_sc_hd__nand3_2 _16469_ (.A(_07338_),
    .B(_07340_),
    .C(_07341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07342_));
 sky130_fd_sc_hd__a21o_2 _16470_ (.A1(_07338_),
    .A2(_07341_),
    .B1(_07340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07343_));
 sky130_fd_sc_hd__a21o_2 _16471_ (.A1(_07338_),
    .A2(_07341_),
    .B1(_07339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07344_));
 sky130_fd_sc_hd__nand2_2 _16472_ (.A(_07338_),
    .B(_07339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07345_));
 sky130_fd_sc_hd__nand3_2 _16473_ (.A(_07338_),
    .B(_07341_),
    .C(_07339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07346_));
 sky130_fd_sc_hd__nand2_2 _16474_ (.A(_07344_),
    .B(_07346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07347_));
 sky130_fd_sc_hd__nand2_2 _16475_ (.A(_07342_),
    .B(_07343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_2 _16476_ (.A(_07256_),
    .B(_07279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_2 _16477_ (.A(_07257_),
    .B(_07349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07350_));
 sky130_fd_sc_hd__a21boi_2 _16478_ (.A1(_07256_),
    .A2(_07279_),
    .B1_N(_07257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07351_));
 sky130_fd_sc_hd__o21a_2 _16479_ (.A1(_07129_),
    .A2(_07262_),
    .B1(_07267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07352_));
 sky130_fd_sc_hd__nand2_2 _16480_ (.A(\a_l[8] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07353_));
 sky130_fd_sc_hd__nand2_2 _16481_ (.A(_07262_),
    .B(_07353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07354_));
 sky130_fd_sc_hd__nand2_2 _16482_ (.A(\a_l[8] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07355_));
 sky130_fd_sc_hd__nand4_2 _16483_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07356_));
 sky130_fd_sc_hd__nand3_2 _16484_ (.A(_07353_),
    .B(\b_h[7] ),
    .C(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07357_));
 sky130_fd_sc_hd__nand3_2 _16485_ (.A(_07262_),
    .B(\b_h[6] ),
    .C(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07358_));
 sky130_fd_sc_hd__o211ai_2 _16486_ (.A1(_09231_),
    .A2(_09613_),
    .B1(_07357_),
    .C1(_07358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07359_));
 sky130_fd_sc_hd__nand4_2 _16487_ (.A(_07354_),
    .B(_07356_),
    .C(\a_l[6] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07360_));
 sky130_fd_sc_hd__o21ai_2 _16488_ (.A1(_07246_),
    .A2(_07242_),
    .B1(_07245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07361_));
 sky130_fd_sc_hd__a21oi_2 _16489_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07362_));
 sky130_fd_sc_hd__a21o_2 _16490_ (.A1(_07359_),
    .A2(_07360_),
    .B1(_07361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07363_));
 sky130_fd_sc_hd__nand3_2 _16491_ (.A(_07361_),
    .B(_07360_),
    .C(_07359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07364_));
 sky130_fd_sc_hd__a21o_2 _16492_ (.A1(_07363_),
    .A2(_07364_),
    .B1(_07352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07365_));
 sky130_fd_sc_hd__nand4_2 _16493_ (.A(_07263_),
    .B(_07267_),
    .C(_07363_),
    .D(_07364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07366_));
 sky130_fd_sc_hd__nand2_2 _16494_ (.A(_07365_),
    .B(_07366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_2 _16495_ (.A1(_07247_),
    .A2(_07250_),
    .B1(_07240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07368_));
 sky130_fd_sc_hd__a32oi_2 _16496_ (.A1(_07227_),
    .A2(_07236_),
    .A3(_07237_),
    .B1(_07251_),
    .B2(_07240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07369_));
 sky130_fd_sc_hd__nand2_2 _16497_ (.A(_07241_),
    .B(_07368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07370_));
 sky130_fd_sc_hd__nor2_2 _16498_ (.A(_09340_),
    .B(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07371_));
 sky130_fd_sc_hd__nand2_2 _16499_ (.A(\a_l[13] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07372_));
 sky130_fd_sc_hd__nand2_2 _16500_ (.A(\a_l[11] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07373_));
 sky130_fd_sc_hd__nand2_2 _16501_ (.A(\a_l[12] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07374_));
 sky130_fd_sc_hd__a22oi_2 _16502_ (.A1(\a_l[12] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_2 _16503_ (.A(_07373_),
    .B(_07374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07376_));
 sky130_fd_sc_hd__nand2_2 _16504_ (.A(\a_l[12] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07377_));
 sky130_fd_sc_hd__nand4_2 _16505_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07378_));
 sky130_fd_sc_hd__nand2_2 _16506_ (.A(_07376_),
    .B(_07378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07379_));
 sky130_fd_sc_hd__o2bb2a_2 _16507_ (.A1_N(_07376_),
    .A2_N(_07378_),
    .B1(_09340_),
    .B2(_09581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07380_));
 sky130_fd_sc_hd__a22o_2 _16508_ (.A1(\a_l[13] ),
    .A2(\b_h[1] ),
    .B1(_07376_),
    .B2(_07378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07381_));
 sky130_fd_sc_hd__o2111ai_2 _16509_ (.A1(_07231_),
    .A2(_07377_),
    .B1(\a_l[13] ),
    .C1(\b_h[1] ),
    .D1(_07376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07382_));
 sky130_fd_sc_hd__nand2_2 _16510_ (.A(_07372_),
    .B(_07378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07383_));
 sky130_fd_sc_hd__nand2_2 _16511_ (.A(_07379_),
    .B(_07371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07384_));
 sky130_fd_sc_hd__a21o_2 _16512_ (.A1(_07229_),
    .A2(_07235_),
    .B1(_07232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07385_));
 sky130_fd_sc_hd__a21oi_2 _16513_ (.A1(_07229_),
    .A2(_07235_),
    .B1(_07232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07386_));
 sky130_fd_sc_hd__o211ai_2 _16514_ (.A1(_07375_),
    .A2(_07383_),
    .B1(_07385_),
    .C1(_07384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07387_));
 sky130_fd_sc_hd__o21ai_2 _16515_ (.A1(_07372_),
    .A2(_07379_),
    .B1(_07386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07388_));
 sky130_fd_sc_hd__nand3_2 _16516_ (.A(_07381_),
    .B(_07382_),
    .C(_07386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07389_));
 sky130_fd_sc_hd__nand2_2 _16517_ (.A(\a_l[9] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07390_));
 sky130_fd_sc_hd__a22oi_2 _16518_ (.A1(\a_l[14] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_2 _16519_ (.A(\a_l[14] ),
    .B(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07392_));
 sky130_fd_sc_hd__and4_2 _16520_ (.A(\a_l[10] ),
    .B(\a_l[14] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07393_));
 sky130_fd_sc_hd__o21a_2 _16521_ (.A1(_06878_),
    .A2(_07392_),
    .B1(_07390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07394_));
 sky130_fd_sc_hd__o21ai_2 _16522_ (.A1(_06878_),
    .A2(_07392_),
    .B1(_07390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07395_));
 sky130_fd_sc_hd__nor2_2 _16523_ (.A(_07391_),
    .B(_07395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07396_));
 sky130_fd_sc_hd__o211a_2 _16524_ (.A1(_07391_),
    .A2(_07393_),
    .B1(\a_l[9] ),
    .C1(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07397_));
 sky130_fd_sc_hd__o21bai_2 _16525_ (.A1(_07391_),
    .A2(_07393_),
    .B1_N(_07390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07398_));
 sky130_fd_sc_hd__o21ai_2 _16526_ (.A1(_07391_),
    .A2(_07395_),
    .B1(_07398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07399_));
 sky130_fd_sc_hd__a21oi_2 _16527_ (.A1(_07387_),
    .A2(_07389_),
    .B1(_07399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07400_));
 sky130_fd_sc_hd__a21o_2 _16528_ (.A1(_07387_),
    .A2(_07389_),
    .B1(_07399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07401_));
 sky130_fd_sc_hd__nand3_2 _16529_ (.A(_07387_),
    .B(_07389_),
    .C(_07399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07402_));
 sky130_fd_sc_hd__o2111ai_2 _16530_ (.A1(_07391_),
    .A2(_07395_),
    .B1(_07398_),
    .C1(_07389_),
    .D1(_07387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07403_));
 sky130_fd_sc_hd__o2bb2ai_2 _16531_ (.A1_N(_07387_),
    .A2_N(_07389_),
    .B1(_07396_),
    .B2(_07397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07404_));
 sky130_fd_sc_hd__nand3_2 _16532_ (.A(_07241_),
    .B(_07368_),
    .C(_07402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07405_));
 sky130_fd_sc_hd__a21oi_2 _16533_ (.A1(_07403_),
    .A2(_07404_),
    .B1(_07370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07406_));
 sky130_fd_sc_hd__nand3_2 _16534_ (.A(_07401_),
    .B(_07402_),
    .C(_07369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07407_));
 sky130_fd_sc_hd__nand3_2 _16535_ (.A(_07370_),
    .B(_07403_),
    .C(_07404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07408_));
 sky130_fd_sc_hd__o21ai_2 _16536_ (.A1(_07400_),
    .A2(_07405_),
    .B1(_07408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07409_));
 sky130_fd_sc_hd__nand2_2 _16537_ (.A(_07408_),
    .B(_07367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07410_));
 sky130_fd_sc_hd__a21o_2 _16538_ (.A1(_07407_),
    .A2(_07408_),
    .B1(_07367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07411_));
 sky130_fd_sc_hd__nand4_2 _16539_ (.A(_07365_),
    .B(_07366_),
    .C(_07407_),
    .D(_07408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07412_));
 sky130_fd_sc_hd__nand2_2 _16540_ (.A(_07409_),
    .B(_07367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07413_));
 sky130_fd_sc_hd__a21oi_2 _16541_ (.A1(_07412_),
    .A2(_07413_),
    .B1(_07350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07414_));
 sky130_fd_sc_hd__o211ai_2 _16542_ (.A1(_07410_),
    .A2(_07406_),
    .B1(_07351_),
    .C1(_07411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07415_));
 sky130_fd_sc_hd__nand3_2 _16543_ (.A(_07350_),
    .B(_07412_),
    .C(_07413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07416_));
 sky130_fd_sc_hd__nand2_2 _16544_ (.A(_07347_),
    .B(_07416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07417_));
 sky130_fd_sc_hd__a22o_2 _16545_ (.A1(_07342_),
    .A2(_07343_),
    .B1(_07415_),
    .B2(_07416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07418_));
 sky130_fd_sc_hd__nand2_2 _16546_ (.A(_07348_),
    .B(_07416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07419_));
 sky130_fd_sc_hd__a22o_2 _16547_ (.A1(_07344_),
    .A2(_07346_),
    .B1(_07415_),
    .B2(_07416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07420_));
 sky130_fd_sc_hd__o211ai_2 _16548_ (.A1(_07417_),
    .A2(_07414_),
    .B1(_07310_),
    .C1(_07418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07421_));
 sky130_fd_sc_hd__a32oi_2 _16549_ (.A1(_07348_),
    .A2(_07415_),
    .A3(_07416_),
    .B1(_07287_),
    .B2(_07285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07422_));
 sky130_fd_sc_hd__o211ai_2 _16550_ (.A1(_07414_),
    .A2(_07419_),
    .B1(_07309_),
    .C1(_07420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07423_));
 sky130_fd_sc_hd__a211oi_2 _16551_ (.A1(_07214_),
    .A2(_07220_),
    .B1(_02589_),
    .C1(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07424_));
 sky130_fd_sc_hd__a22o_2 _16552_ (.A1(_02588_),
    .A2(_06401_),
    .B1(_07219_),
    .B2(_07212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07425_));
 sky130_fd_sc_hd__o21ba_2 _16553_ (.A1(_07213_),
    .A2(_07425_),
    .B1_N(_07424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07426_));
 sky130_fd_sc_hd__o21bai_2 _16554_ (.A1(_07213_),
    .A2(_07425_),
    .B1_N(_07424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07427_));
 sky130_fd_sc_hd__a21oi_2 _16555_ (.A1(_07421_),
    .A2(_07423_),
    .B1(_07427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07428_));
 sky130_fd_sc_hd__and3_2 _16556_ (.A(_07421_),
    .B(_07423_),
    .C(_07427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07429_));
 sky130_fd_sc_hd__nand3_2 _16557_ (.A(_07421_),
    .B(_07423_),
    .C(_07427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07430_));
 sky130_fd_sc_hd__a21boi_2 _16558_ (.A1(_07292_),
    .A2(_07294_),
    .B1_N(_07289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07431_));
 sky130_fd_sc_hd__nand3b_2 _16559_ (.A_N(_07428_),
    .B(_07430_),
    .C(_07431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07432_));
 sky130_fd_sc_hd__o21bai_2 _16560_ (.A1(_07428_),
    .A2(_07429_),
    .B1_N(_07431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07433_));
 sky130_fd_sc_hd__nand3_2 _16561_ (.A(_07302_),
    .B(_07432_),
    .C(_07433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07434_));
 sky130_fd_sc_hd__a32o_2 _16562_ (.A1(_07297_),
    .A2(_07299_),
    .A3(_07298_),
    .B1(_07433_),
    .B2(_07432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07435_));
 sky130_fd_sc_hd__a211oi_2 _16563_ (.A1(_07051_),
    .A2(_07177_),
    .B1(_07178_),
    .C1(_07304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07436_));
 sky130_fd_sc_hd__o2111a_2 _16564_ (.A1(_07302_),
    .A2(_07305_),
    .B1(_07306_),
    .C1(_07182_),
    .D1(_07181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07437_));
 sky130_fd_sc_hd__nand2_2 _16565_ (.A(_07060_),
    .B(_07437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07438_));
 sky130_fd_sc_hd__a21o_2 _16566_ (.A1(_07060_),
    .A2(_07437_),
    .B1(_07436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07439_));
 sky130_fd_sc_hd__a221o_2 _16567_ (.A1(_07434_),
    .A2(_07435_),
    .B1(_07184_),
    .B2(_07307_),
    .C1(_07436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07440_));
 sky130_fd_sc_hd__nand3_2 _16568_ (.A(_07434_),
    .B(_07435_),
    .C(_07439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07441_));
 sky130_fd_sc_hd__and3_2 _16569_ (.A(_09690_),
    .B(_07440_),
    .C(_07441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00352_));
 sky130_fd_sc_hd__a22o_2 _16570_ (.A1(_07420_),
    .A2(_07422_),
    .B1(_07421_),
    .B2(_07426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07442_));
 sky130_fd_sc_hd__a22oi_2 _16571_ (.A1(_07420_),
    .A2(_07422_),
    .B1(_07421_),
    .B2(_07426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07443_));
 sky130_fd_sc_hd__a2bb2o_2 _16572_ (.A1_N(_07315_),
    .A2_N(_07316_),
    .B1(_07341_),
    .B2(_07345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07444_));
 sky130_fd_sc_hd__o2111ai_2 _16573_ (.A1(_02589_),
    .A2(_06441_),
    .B1(_07317_),
    .C1(_07341_),
    .D1(_07345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_2 _16574_ (.A(_07444_),
    .B(_07445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07446_));
 sky130_fd_sc_hd__nand2_2 _16575_ (.A(\a_l[0] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07447_));
 sky130_fd_sc_hd__a21o_2 _16576_ (.A1(_07444_),
    .A2(_07445_),
    .B1(_07447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07448_));
 sky130_fd_sc_hd__o211ai_2 _16577_ (.A1(_09166_),
    .A2(_09679_),
    .B1(_07444_),
    .C1(_07445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07449_));
 sky130_fd_sc_hd__nand2_2 _16578_ (.A(_07448_),
    .B(_07449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07450_));
 sky130_fd_sc_hd__a21oi_2 _16579_ (.A1(_07348_),
    .A2(_07416_),
    .B1(_07414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07451_));
 sky130_fd_sc_hd__a21o_2 _16580_ (.A1(_07348_),
    .A2(_07416_),
    .B1(_07414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07452_));
 sky130_fd_sc_hd__o21ai_2 _16581_ (.A1(_07352_),
    .A2(_07362_),
    .B1(_07364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07453_));
 sky130_fd_sc_hd__o21a_2 _16582_ (.A1(_07352_),
    .A2(_07362_),
    .B1(_07364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07454_));
 sky130_fd_sc_hd__nand2_2 _16583_ (.A(\a_l[4] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07455_));
 sky130_fd_sc_hd__nand2_2 _16584_ (.A(\a_l[5] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07456_));
 sky130_fd_sc_hd__nand2_2 _16585_ (.A(\a_l[6] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07457_));
 sky130_fd_sc_hd__a22oi_2 _16586_ (.A1(\a_l[6] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07458_));
 sky130_fd_sc_hd__nand2_2 _16587_ (.A(_07456_),
    .B(_07457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07459_));
 sky130_fd_sc_hd__nand4_2 _16588_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07460_));
 sky130_fd_sc_hd__a22o_2 _16589_ (.A1(\a_l[4] ),
    .A2(\b_h[11] ),
    .B1(_07459_),
    .B2(_07460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07461_));
 sky130_fd_sc_hd__nand4_2 _16590_ (.A(_07459_),
    .B(_07460_),
    .C(\a_l[4] ),
    .D(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07462_));
 sky130_fd_sc_hd__a21o_2 _16591_ (.A1(_07459_),
    .A2(_07460_),
    .B1(_07455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07463_));
 sky130_fd_sc_hd__o211ai_2 _16592_ (.A1(_09199_),
    .A2(_09646_),
    .B1(_07459_),
    .C1(_07460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07464_));
 sky130_fd_sc_hd__o2bb2ai_2 _16593_ (.A1_N(_07327_),
    .A2_N(_07324_),
    .B1(_09624_),
    .B2(_07325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07465_));
 sky130_fd_sc_hd__a21boi_2 _16594_ (.A1(_07324_),
    .A2(_07327_),
    .B1_N(_07326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07466_));
 sky130_fd_sc_hd__and3_2 _16595_ (.A(_07463_),
    .B(_07464_),
    .C(_07466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07467_));
 sky130_fd_sc_hd__nand3_2 _16596_ (.A(_07463_),
    .B(_07464_),
    .C(_07466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07468_));
 sky130_fd_sc_hd__nand3_2 _16597_ (.A(_07461_),
    .B(_07462_),
    .C(_07465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07469_));
 sky130_fd_sc_hd__nand2_2 _16598_ (.A(_07468_),
    .B(_07469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07470_));
 sky130_fd_sc_hd__a22oi_2 _16599_ (.A1(\a_l[3] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07471_));
 sky130_fd_sc_hd__and4_2 _16600_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07472_));
 sky130_fd_sc_hd__nand4_2 _16601_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07473_));
 sky130_fd_sc_hd__nand4b_2 _16602_ (.A_N(_07471_),
    .B(_07473_),
    .C(\a_l[1] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07474_));
 sky130_fd_sc_hd__o2bb2ai_2 _16603_ (.A1_N(\a_l[1] ),
    .A2_N(\b_h[14] ),
    .B1(_07471_),
    .B2(_07472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07475_));
 sky130_fd_sc_hd__a211oi_2 _16604_ (.A1(\a_l[1] ),
    .A2(\b_h[14] ),
    .B1(_07471_),
    .C1(_07472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07476_));
 sky130_fd_sc_hd__o211a_2 _16605_ (.A1(_07471_),
    .A2(_07472_),
    .B1(\a_l[1] ),
    .C1(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07477_));
 sky130_fd_sc_hd__nand2_2 _16606_ (.A(_07474_),
    .B(_07475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07478_));
 sky130_fd_sc_hd__o2bb2ai_2 _16607_ (.A1_N(_07468_),
    .A2_N(_07469_),
    .B1(_07476_),
    .B2(_07477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07479_));
 sky130_fd_sc_hd__nand3_2 _16608_ (.A(_07468_),
    .B(_07469_),
    .C(_07478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07480_));
 sky130_fd_sc_hd__nand4_2 _16609_ (.A(_07468_),
    .B(_07469_),
    .C(_07474_),
    .D(_07475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07481_));
 sky130_fd_sc_hd__nand2_2 _16610_ (.A(_07470_),
    .B(_07478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07482_));
 sky130_fd_sc_hd__nand3_2 _16611_ (.A(_07482_),
    .B(_07453_),
    .C(_07481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07483_));
 sky130_fd_sc_hd__nand3_2 _16612_ (.A(_07454_),
    .B(_07479_),
    .C(_07480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07484_));
 sky130_fd_sc_hd__o21ai_2 _16613_ (.A1(_07332_),
    .A2(_07320_),
    .B1(_07331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07485_));
 sky130_fd_sc_hd__a21o_2 _16614_ (.A1(_07483_),
    .A2(_07484_),
    .B1(_07485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07486_));
 sky130_fd_sc_hd__nand2_2 _16615_ (.A(_07484_),
    .B(_07485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07487_));
 sky130_fd_sc_hd__nand3_2 _16616_ (.A(_07483_),
    .B(_07484_),
    .C(_07485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07488_));
 sky130_fd_sc_hd__nand2_2 _16617_ (.A(_07486_),
    .B(_07488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07489_));
 sky130_fd_sc_hd__o2bb2ai_2 _16618_ (.A1_N(_07367_),
    .A2_N(_07408_),
    .B1(_07405_),
    .B2(_07400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07490_));
 sky130_fd_sc_hd__a21oi_2 _16619_ (.A1(_07367_),
    .A2(_07408_),
    .B1(_07406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07491_));
 sky130_fd_sc_hd__o21ai_2 _16620_ (.A1(_07260_),
    .A2(_07355_),
    .B1(_07360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07492_));
 sky130_fd_sc_hd__nor2_2 _16621_ (.A(_07390_),
    .B(_07391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07493_));
 sky130_fd_sc_hd__nand2_2 _16622_ (.A(\a_l[7] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07494_));
 sky130_fd_sc_hd__nand2_2 _16623_ (.A(\a_l[9] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07495_));
 sky130_fd_sc_hd__a22oi_2 _16624_ (.A1(\a_l[9] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07496_));
 sky130_fd_sc_hd__nand2_2 _16625_ (.A(_07355_),
    .B(_07495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07497_));
 sky130_fd_sc_hd__nand2_2 _16626_ (.A(\a_l[9] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07498_));
 sky130_fd_sc_hd__nand4_2 _16627_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07499_));
 sky130_fd_sc_hd__o2111ai_2 _16628_ (.A1(_07353_),
    .A2(_07498_),
    .B1(\a_l[7] ),
    .C1(\b_h[8] ),
    .D1(_07497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07500_));
 sky130_fd_sc_hd__a22o_2 _16629_ (.A1(\a_l[7] ),
    .A2(\b_h[8] ),
    .B1(_07497_),
    .B2(_07499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07501_));
 sky130_fd_sc_hd__nand3_2 _16630_ (.A(_07395_),
    .B(_07500_),
    .C(_07501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07502_));
 sky130_fd_sc_hd__o211ai_2 _16631_ (.A1(_07393_),
    .A2(_07493_),
    .B1(_07500_),
    .C1(_07501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07503_));
 sky130_fd_sc_hd__o221ai_2 _16632_ (.A1(_09242_),
    .A2(_09613_),
    .B1(_07353_),
    .B2(_07498_),
    .C1(_07497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07504_));
 sky130_fd_sc_hd__a21o_2 _16633_ (.A1(_07497_),
    .A2(_07499_),
    .B1(_07494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07505_));
 sky130_fd_sc_hd__o211ai_2 _16634_ (.A1(_07391_),
    .A2(_07394_),
    .B1(_07504_),
    .C1(_07505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07506_));
 sky130_fd_sc_hd__a21o_2 _16635_ (.A1(_07503_),
    .A2(_07506_),
    .B1(_07492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07507_));
 sky130_fd_sc_hd__o211ai_2 _16636_ (.A1(_07391_),
    .A2(_07502_),
    .B1(_07506_),
    .C1(_07492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07508_));
 sky130_fd_sc_hd__nand2_2 _16637_ (.A(_07507_),
    .B(_07508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07509_));
 sky130_fd_sc_hd__o2bb2ai_2 _16638_ (.A1_N(_07399_),
    .A2_N(_07387_),
    .B1(_07380_),
    .B2(_07388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07510_));
 sky130_fd_sc_hd__a21boi_2 _16639_ (.A1(_07387_),
    .A2(_07399_),
    .B1_N(_07389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07511_));
 sky130_fd_sc_hd__nand2_2 _16640_ (.A(\a_l[10] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07512_));
 sky130_fd_sc_hd__nand2_2 _16641_ (.A(\a_l[15] ),
    .B(\b_h[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07513_));
 sky130_fd_sc_hd__a22oi_2 _16642_ (.A1(\a_l[15] ),
    .A2(\b_h[0] ),
    .B1(\b_h[4] ),
    .B2(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07514_));
 sky130_fd_sc_hd__nand2_2 _16643_ (.A(_06999_),
    .B(_07513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07515_));
 sky130_fd_sc_hd__nand4_2 _16644_ (.A(\a_l[11] ),
    .B(\a_l[15] ),
    .C(\b_h[0] ),
    .D(\b_h[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07516_));
 sky130_fd_sc_hd__a21o_2 _16645_ (.A1(_07515_),
    .A2(_07516_),
    .B1(_07512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07517_));
 sky130_fd_sc_hd__o21ai_2 _16646_ (.A1(_06999_),
    .A2(_07513_),
    .B1(_07512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07518_));
 sky130_fd_sc_hd__o21ai_2 _16647_ (.A1(_07514_),
    .A2(_07518_),
    .B1(_07517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07519_));
 sky130_fd_sc_hd__o21a_2 _16648_ (.A1(_07514_),
    .A2(_07518_),
    .B1(_07517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07520_));
 sky130_fd_sc_hd__nand2_2 _16649_ (.A(_07376_),
    .B(_07383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07521_));
 sky130_fd_sc_hd__a21oi_2 _16650_ (.A1(_07372_),
    .A2(_07378_),
    .B1(_07375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07522_));
 sky130_fd_sc_hd__and2_2 _16651_ (.A(\a_l[14] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07523_));
 sky130_fd_sc_hd__nand2_2 _16652_ (.A(\a_l[14] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07524_));
 sky130_fd_sc_hd__nand2_2 _16653_ (.A(\a_l[13] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07525_));
 sky130_fd_sc_hd__a22oi_2 _16654_ (.A1(\a_l[13] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07526_));
 sky130_fd_sc_hd__nand2_2 _16655_ (.A(_07377_),
    .B(_07525_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07527_));
 sky130_fd_sc_hd__nand4_2 _16656_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07528_));
 sky130_fd_sc_hd__nand2_2 _16657_ (.A(_07527_),
    .B(_07528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07529_));
 sky130_fd_sc_hd__a21oi_2 _16658_ (.A1(_07527_),
    .A2(_07528_),
    .B1(_07523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07530_));
 sky130_fd_sc_hd__a22o_2 _16659_ (.A1(\a_l[14] ),
    .A2(\b_h[1] ),
    .B1(_07527_),
    .B2(_07528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07531_));
 sky130_fd_sc_hd__nand4_2 _16660_ (.A(_07527_),
    .B(_07528_),
    .C(\a_l[14] ),
    .D(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07532_));
 sky130_fd_sc_hd__nand2_2 _16661_ (.A(_07529_),
    .B(_07523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07533_));
 sky130_fd_sc_hd__nand2_2 _16662_ (.A(_07524_),
    .B(_07528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07534_));
 sky130_fd_sc_hd__nand3_2 _16663_ (.A(_07524_),
    .B(_07527_),
    .C(_07528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07535_));
 sky130_fd_sc_hd__nand2_2 _16664_ (.A(_07522_),
    .B(_07532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07536_));
 sky130_fd_sc_hd__and3_2 _16665_ (.A(_07533_),
    .B(_07535_),
    .C(_07521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07537_));
 sky130_fd_sc_hd__nand3_2 _16666_ (.A(_07533_),
    .B(_07535_),
    .C(_07521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07538_));
 sky130_fd_sc_hd__o21ai_2 _16667_ (.A1(_07530_),
    .A2(_07536_),
    .B1(_07538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_2 _16668_ (.A(_07520_),
    .B(_07539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07540_));
 sky130_fd_sc_hd__o211ai_2 _16669_ (.A1(_07530_),
    .A2(_07536_),
    .B1(_07519_),
    .C1(_07538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07541_));
 sky130_fd_sc_hd__o211ai_2 _16670_ (.A1(_07530_),
    .A2(_07536_),
    .B1(_07538_),
    .C1(_07520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07542_));
 sky130_fd_sc_hd__nand2_2 _16671_ (.A(_07539_),
    .B(_07519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07543_));
 sky130_fd_sc_hd__a21oi_2 _16672_ (.A1(_07519_),
    .A2(_07539_),
    .B1(_07510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07544_));
 sky130_fd_sc_hd__and3_2 _16673_ (.A(_07511_),
    .B(_07542_),
    .C(_07543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07545_));
 sky130_fd_sc_hd__nand3_2 _16674_ (.A(_07511_),
    .B(_07542_),
    .C(_07543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07546_));
 sky130_fd_sc_hd__nand3_2 _16675_ (.A(_07540_),
    .B(_07541_),
    .C(_07510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07547_));
 sky130_fd_sc_hd__a32oi_2 _16676_ (.A1(_07540_),
    .A2(_07541_),
    .A3(_07510_),
    .B1(_07508_),
    .B2(_07507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07548_));
 sky130_fd_sc_hd__nand3_2 _16677_ (.A(_07509_),
    .B(_07546_),
    .C(_07547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07549_));
 sky130_fd_sc_hd__inv_2 _16678_ (.A(_07549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07550_));
 sky130_fd_sc_hd__a21o_2 _16679_ (.A1(_07546_),
    .A2(_07547_),
    .B1(_07509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07551_));
 sky130_fd_sc_hd__a22o_2 _16680_ (.A1(_07507_),
    .A2(_07508_),
    .B1(_07546_),
    .B2(_07547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07552_));
 sky130_fd_sc_hd__nand4_2 _16681_ (.A(_07507_),
    .B(_07508_),
    .C(_07546_),
    .D(_07547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07553_));
 sky130_fd_sc_hd__nand2_2 _16682_ (.A(_07491_),
    .B(_07551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07554_));
 sky130_fd_sc_hd__nand3_2 _16683_ (.A(_07491_),
    .B(_07549_),
    .C(_07551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07555_));
 sky130_fd_sc_hd__and3_2 _16684_ (.A(_07552_),
    .B(_07553_),
    .C(_07490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07556_));
 sky130_fd_sc_hd__nand3_2 _16685_ (.A(_07552_),
    .B(_07553_),
    .C(_07490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07557_));
 sky130_fd_sc_hd__o211ai_2 _16686_ (.A1(_07550_),
    .A2(_07554_),
    .B1(_07557_),
    .C1(_07489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07558_));
 sky130_fd_sc_hd__a21o_2 _16687_ (.A1(_07555_),
    .A2(_07557_),
    .B1(_07489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07559_));
 sky130_fd_sc_hd__and4_2 _16688_ (.A(_07486_),
    .B(_07488_),
    .C(_07555_),
    .D(_07557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07560_));
 sky130_fd_sc_hd__nand4_2 _16689_ (.A(_07486_),
    .B(_07488_),
    .C(_07555_),
    .D(_07557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07561_));
 sky130_fd_sc_hd__a22o_2 _16690_ (.A1(_07486_),
    .A2(_07488_),
    .B1(_07555_),
    .B2(_07557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07562_));
 sky130_fd_sc_hd__nand2_2 _16691_ (.A(_07452_),
    .B(_07562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07563_));
 sky130_fd_sc_hd__nand3_2 _16692_ (.A(_07452_),
    .B(_07561_),
    .C(_07562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07564_));
 sky130_fd_sc_hd__nand3_2 _16693_ (.A(_07559_),
    .B(_07451_),
    .C(_07558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07565_));
 sky130_fd_sc_hd__nand2_2 _16694_ (.A(_07564_),
    .B(_07565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07566_));
 sky130_fd_sc_hd__nand2_2 _16695_ (.A(_07566_),
    .B(_07450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07567_));
 sky130_fd_sc_hd__nand3b_2 _16696_ (.A_N(_07450_),
    .B(_07564_),
    .C(_07565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07568_));
 sky130_fd_sc_hd__and3_2 _16697_ (.A(_07564_),
    .B(_07565_),
    .C(_07450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07569_));
 sky130_fd_sc_hd__o211ai_2 _16698_ (.A1(_07560_),
    .A2(_07563_),
    .B1(_07565_),
    .C1(_07450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07570_));
 sky130_fd_sc_hd__a21o_2 _16699_ (.A1(_07564_),
    .A2(_07565_),
    .B1(_07450_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07571_));
 sky130_fd_sc_hd__nand2_2 _16700_ (.A(_07442_),
    .B(_07571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07572_));
 sky130_fd_sc_hd__nand3_2 _16701_ (.A(_07442_),
    .B(_07570_),
    .C(_07571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07573_));
 sky130_fd_sc_hd__nand3_2 _16702_ (.A(_07443_),
    .B(_07567_),
    .C(_07568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07574_));
 sky130_fd_sc_hd__a21bo_2 _16703_ (.A1(_07573_),
    .A2(_07574_),
    .B1_N(_07424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07575_));
 sky130_fd_sc_hd__nand3b_2 _16704_ (.A_N(_07424_),
    .B(_07573_),
    .C(_07574_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07576_));
 sky130_fd_sc_hd__nand2_2 _16705_ (.A(_07575_),
    .B(_07576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07577_));
 sky130_fd_sc_hd__nand3_2 _16706_ (.A(_07433_),
    .B(_07575_),
    .C(_07576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07578_));
 sky130_fd_sc_hd__a32oi_2 _16707_ (.A1(_07433_),
    .A2(_07575_),
    .A3(_07576_),
    .B1(_07434_),
    .B2(_07441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07579_));
 sky130_fd_sc_hd__a21o_2 _16708_ (.A1(_07575_),
    .A2(_07576_),
    .B1(_07433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07580_));
 sky130_fd_sc_hd__nand2_2 _16709_ (.A(_07578_),
    .B(_07580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07581_));
 sky130_fd_sc_hd__a311oi_2 _16710_ (.A1(_07434_),
    .A2(_07441_),
    .A3(_07581_),
    .B1(_07579_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_2 _16711_ (.A(_07433_),
    .B(_07434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07582_));
 sky130_fd_sc_hd__a21oi_2 _16712_ (.A1(_07577_),
    .A2(_07582_),
    .B1(_07436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07583_));
 sky130_fd_sc_hd__nand2_2 _16713_ (.A(_07438_),
    .B(_07583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07584_));
 sky130_fd_sc_hd__nand2_2 _16714_ (.A(_07435_),
    .B(_07578_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07585_));
 sky130_fd_sc_hd__nand2_2 _16715_ (.A(_07580_),
    .B(_07585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07586_));
 sky130_fd_sc_hd__a22oi_2 _16716_ (.A1(_07580_),
    .A2(_07585_),
    .B1(_07438_),
    .B2(_07583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07587_));
 sky130_fd_sc_hd__o2bb2ai_2 _16717_ (.A1_N(_07450_),
    .A2_N(_07565_),
    .B1(_07560_),
    .B2(_07563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07588_));
 sky130_fd_sc_hd__a21boi_2 _16718_ (.A1(_07450_),
    .A2(_07565_),
    .B1_N(_07564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07589_));
 sky130_fd_sc_hd__a31oi_2 _16719_ (.A1(_07491_),
    .A2(_07549_),
    .A3(_07551_),
    .B1(_07489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07590_));
 sky130_fd_sc_hd__o2bb2ai_2 _16720_ (.A1_N(_07489_),
    .A2_N(_07557_),
    .B1(_07554_),
    .B2(_07550_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07591_));
 sky130_fd_sc_hd__o2bb2ai_2 _16721_ (.A1_N(_07492_),
    .A2_N(_07506_),
    .B1(_07391_),
    .B2(_07502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07592_));
 sky130_fd_sc_hd__a22o_2 _16722_ (.A1(\a_l[4] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07593_));
 sky130_fd_sc_hd__and4_2 _16723_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07594_));
 sky130_fd_sc_hd__nand4_2 _16724_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07595_));
 sky130_fd_sc_hd__nand2_2 _16725_ (.A(\a_l[2] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07596_));
 sky130_fd_sc_hd__o211ai_2 _16726_ (.A1(_09144_),
    .A2(_09668_),
    .B1(_07593_),
    .C1(_07595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07597_));
 sky130_fd_sc_hd__a21o_2 _16727_ (.A1(_07593_),
    .A2(_07595_),
    .B1(_07596_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07598_));
 sky130_fd_sc_hd__nand2_2 _16728_ (.A(_07597_),
    .B(_07598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07599_));
 sky130_fd_sc_hd__o21ai_2 _16729_ (.A1(_07455_),
    .A2(_07458_),
    .B1(_07460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07600_));
 sky130_fd_sc_hd__o21a_2 _16730_ (.A1(_07455_),
    .A2(_07458_),
    .B1(_07460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07601_));
 sky130_fd_sc_hd__nor2_2 _16731_ (.A(_09210_),
    .B(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07602_));
 sky130_fd_sc_hd__nand2_2 _16732_ (.A(\a_l[5] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07603_));
 sky130_fd_sc_hd__nand2_2 _16733_ (.A(\a_l[6] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07604_));
 sky130_fd_sc_hd__nand2_2 _16734_ (.A(\a_l[7] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07605_));
 sky130_fd_sc_hd__nand4_2 _16735_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07606_));
 sky130_fd_sc_hd__a22oi_2 _16736_ (.A1(\a_l[7] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07607_));
 sky130_fd_sc_hd__nand2_2 _16737_ (.A(_07604_),
    .B(_07605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07608_));
 sky130_fd_sc_hd__o21ai_2 _16738_ (.A1(_02338_),
    .A2(_06761_),
    .B1(_07608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07609_));
 sky130_fd_sc_hd__o21ai_2 _16739_ (.A1(_09210_),
    .A2(_09646_),
    .B1(_07609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07610_));
 sky130_fd_sc_hd__o2111ai_2 _16740_ (.A1(_02338_),
    .A2(_06761_),
    .B1(\a_l[5] ),
    .C1(\b_h[11] ),
    .D1(_07608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07611_));
 sky130_fd_sc_hd__nand2_2 _16741_ (.A(_07609_),
    .B(_07602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07612_));
 sky130_fd_sc_hd__o221ai_2 _16742_ (.A1(_09210_),
    .A2(_09646_),
    .B1(_02338_),
    .B2(_06761_),
    .C1(_07608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07613_));
 sky130_fd_sc_hd__nand3_2 _16743_ (.A(_07601_),
    .B(_07612_),
    .C(_07613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07614_));
 sky130_fd_sc_hd__nand3_2 _16744_ (.A(_07610_),
    .B(_07611_),
    .C(_07600_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07615_));
 sky130_fd_sc_hd__nand3_2 _16745_ (.A(_07599_),
    .B(_07614_),
    .C(_07615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07616_));
 sky130_fd_sc_hd__a21o_2 _16746_ (.A1(_07614_),
    .A2(_07615_),
    .B1(_07599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07617_));
 sky130_fd_sc_hd__a22o_2 _16747_ (.A1(_07597_),
    .A2(_07598_),
    .B1(_07614_),
    .B2(_07615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07618_));
 sky130_fd_sc_hd__nand4_2 _16748_ (.A(_07597_),
    .B(_07598_),
    .C(_07614_),
    .D(_07615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07619_));
 sky130_fd_sc_hd__nand3_2 _16749_ (.A(_07617_),
    .B(_07592_),
    .C(_07616_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07620_));
 sky130_fd_sc_hd__nand3b_2 _16750_ (.A_N(_07592_),
    .B(_07618_),
    .C(_07619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07621_));
 sky130_fd_sc_hd__o21a_2 _16751_ (.A1(_07478_),
    .A2(_07467_),
    .B1(_07469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07622_));
 sky130_fd_sc_hd__o21ai_2 _16752_ (.A1(_07478_),
    .A2(_07467_),
    .B1(_07469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07623_));
 sky130_fd_sc_hd__a21oi_2 _16753_ (.A1(_07620_),
    .A2(_07621_),
    .B1(_07622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07624_));
 sky130_fd_sc_hd__and3_2 _16754_ (.A(_07620_),
    .B(_07621_),
    .C(_07622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07625_));
 sky130_fd_sc_hd__a21o_2 _16755_ (.A1(_07620_),
    .A2(_07621_),
    .B1(_07623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07626_));
 sky130_fd_sc_hd__nand3_2 _16756_ (.A(_07620_),
    .B(_07621_),
    .C(_07623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07627_));
 sky130_fd_sc_hd__nand2_2 _16757_ (.A(_07626_),
    .B(_07627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07628_));
 sky130_fd_sc_hd__a22oi_2 _16758_ (.A1(_07544_),
    .A2(_07542_),
    .B1(_07509_),
    .B2(_07547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07629_));
 sky130_fd_sc_hd__a31oi_2 _16759_ (.A1(_07522_),
    .A2(_07531_),
    .A3(_07532_),
    .B1(_07519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07630_));
 sky130_fd_sc_hd__o2bb2ai_2 _16760_ (.A1_N(_07519_),
    .A2_N(_07538_),
    .B1(_07536_),
    .B2(_07530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_2 _16761_ (.A(\a_l[12] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07632_));
 sky130_fd_sc_hd__and4_2 _16762_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07633_));
 sky130_fd_sc_hd__or2_2 _16763_ (.A(_06999_),
    .B(_07632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07634_));
 sky130_fd_sc_hd__a22oi_2 _16764_ (.A1(\a_l[12] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07635_));
 sky130_fd_sc_hd__nor2_2 _16765_ (.A(_07633_),
    .B(_07635_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07636_));
 sky130_fd_sc_hd__o21ai_2 _16766_ (.A1(_07524_),
    .A2(_07526_),
    .B1(_07528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_2 _16767_ (.A(_07527_),
    .B(_07534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07638_));
 sky130_fd_sc_hd__and2_2 _16768_ (.A(\a_l[15] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07639_));
 sky130_fd_sc_hd__nand2_2 _16769_ (.A(\a_l[15] ),
    .B(\b_h[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07640_));
 sky130_fd_sc_hd__nand2_2 _16770_ (.A(\a_l[13] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07641_));
 sky130_fd_sc_hd__nand2_2 _16771_ (.A(\a_l[14] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07642_));
 sky130_fd_sc_hd__a22oi_2 _16772_ (.A1(\a_l[14] ),
    .A2(\b_h[2] ),
    .B1(\b_h[3] ),
    .B2(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07643_));
 sky130_fd_sc_hd__nand2_2 _16773_ (.A(_07641_),
    .B(_07642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07644_));
 sky130_fd_sc_hd__nand2_2 _16774_ (.A(\a_l[14] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07645_));
 sky130_fd_sc_hd__and4_2 _16775_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07646_));
 sky130_fd_sc_hd__nand4_2 _16776_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07647_));
 sky130_fd_sc_hd__a21oi_2 _16777_ (.A1(_07644_),
    .A2(_07647_),
    .B1(_07639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07648_));
 sky130_fd_sc_hd__a21o_2 _16778_ (.A1(_07644_),
    .A2(_07647_),
    .B1(_07639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07649_));
 sky130_fd_sc_hd__nand3_2 _16779_ (.A(_07644_),
    .B(_07647_),
    .C(_07639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07650_));
 sky130_fd_sc_hd__a21o_2 _16780_ (.A1(_07644_),
    .A2(_07647_),
    .B1(_07640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07651_));
 sky130_fd_sc_hd__o21a_2 _16781_ (.A1(_07641_),
    .A2(_07642_),
    .B1(_07640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07652_));
 sky130_fd_sc_hd__nand2_2 _16782_ (.A(_07640_),
    .B(_07647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07653_));
 sky130_fd_sc_hd__nand3_2 _16783_ (.A(_07527_),
    .B(_07534_),
    .C(_07650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07654_));
 sky130_fd_sc_hd__nand3_2 _16784_ (.A(_07649_),
    .B(_07650_),
    .C(_07637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07655_));
 sky130_fd_sc_hd__o211ai_2 _16785_ (.A1(_07653_),
    .A2(_07643_),
    .B1(_07638_),
    .C1(_07651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07656_));
 sky130_fd_sc_hd__o21ai_2 _16786_ (.A1(_07648_),
    .A2(_07654_),
    .B1(_07656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07657_));
 sky130_fd_sc_hd__nand2_2 _16787_ (.A(_07656_),
    .B(_07636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07658_));
 sky130_fd_sc_hd__o211a_2 _16788_ (.A1(_07648_),
    .A2(_07654_),
    .B1(_07636_),
    .C1(_07656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07659_));
 sky130_fd_sc_hd__o211ai_2 _16789_ (.A1(_07648_),
    .A2(_07654_),
    .B1(_07636_),
    .C1(_07656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07660_));
 sky130_fd_sc_hd__a21oi_2 _16790_ (.A1(_07655_),
    .A2(_07656_),
    .B1(_07636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07661_));
 sky130_fd_sc_hd__o21ai_2 _16791_ (.A1(_07633_),
    .A2(_07635_),
    .B1(_07657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07662_));
 sky130_fd_sc_hd__nor2_2 _16792_ (.A(_07659_),
    .B(_07661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07663_));
 sky130_fd_sc_hd__nand3_2 _16793_ (.A(_07662_),
    .B(_07631_),
    .C(_07660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07664_));
 sky130_fd_sc_hd__o22ai_2 _16794_ (.A1(_07537_),
    .A2(_07630_),
    .B1(_07659_),
    .B2(_07661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07665_));
 sky130_fd_sc_hd__a21oi_2 _16795_ (.A1(_07512_),
    .A2(_07516_),
    .B1(_07514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07666_));
 sky130_fd_sc_hd__nand2_2 _16796_ (.A(\a_l[8] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07667_));
 sky130_fd_sc_hd__nand2_2 _16797_ (.A(\a_l[10] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07668_));
 sky130_fd_sc_hd__a22oi_2 _16798_ (.A1(\a_l[10] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07669_));
 sky130_fd_sc_hd__nand2_2 _16799_ (.A(_07498_),
    .B(_07668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07670_));
 sky130_fd_sc_hd__nand2_2 _16800_ (.A(\a_l[10] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07671_));
 sky130_fd_sc_hd__nand4_2 _16801_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07672_));
 sky130_fd_sc_hd__o2bb2ai_2 _16802_ (.A1_N(_07670_),
    .A2_N(_07672_),
    .B1(_09253_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07673_));
 sky130_fd_sc_hd__and4_2 _16803_ (.A(_07670_),
    .B(_07672_),
    .C(\a_l[8] ),
    .D(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07674_));
 sky130_fd_sc_hd__o2111ai_2 _16804_ (.A1(_07495_),
    .A2(_07671_),
    .B1(\a_l[8] ),
    .C1(\b_h[8] ),
    .D1(_07670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07675_));
 sky130_fd_sc_hd__o221ai_2 _16805_ (.A1(_09253_),
    .A2(_09613_),
    .B1(_07495_),
    .B2(_07671_),
    .C1(_07670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07676_));
 sky130_fd_sc_hd__a21o_2 _16806_ (.A1(_07670_),
    .A2(_07672_),
    .B1(_07667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07677_));
 sky130_fd_sc_hd__nand3b_2 _16807_ (.A_N(_07666_),
    .B(_07676_),
    .C(_07677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_2 _16808_ (.A(_07666_),
    .B(_07673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07679_));
 sky130_fd_sc_hd__and3_2 _16809_ (.A(_07666_),
    .B(_07673_),
    .C(_07675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07680_));
 sky130_fd_sc_hd__nand3_2 _16810_ (.A(_07666_),
    .B(_07673_),
    .C(_07675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07681_));
 sky130_fd_sc_hd__o22a_2 _16811_ (.A1(_09242_),
    .A2(_09613_),
    .B1(_07353_),
    .B2(_07498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07682_));
 sky130_fd_sc_hd__a21oi_2 _16812_ (.A1(_07494_),
    .A2(_07499_),
    .B1(_07496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07683_));
 sky130_fd_sc_hd__o2bb2a_2 _16813_ (.A1_N(_07678_),
    .A2_N(_07681_),
    .B1(_07682_),
    .B2(_07496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07684_));
 sky130_fd_sc_hd__o2bb2ai_2 _16814_ (.A1_N(_07678_),
    .A2_N(_07681_),
    .B1(_07682_),
    .B2(_07496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07685_));
 sky130_fd_sc_hd__nand2_2 _16815_ (.A(_07678_),
    .B(_07683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07686_));
 sky130_fd_sc_hd__and3_2 _16816_ (.A(_07678_),
    .B(_07681_),
    .C(_07683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07687_));
 sky130_fd_sc_hd__a221oi_2 _16817_ (.A1(_07494_),
    .A2(_07499_),
    .B1(_07678_),
    .B2(_07681_),
    .C1(_07496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07688_));
 sky130_fd_sc_hd__o211a_2 _16818_ (.A1(_07496_),
    .A2(_07682_),
    .B1(_07681_),
    .C1(_07678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07689_));
 sky130_fd_sc_hd__o21ai_2 _16819_ (.A1(_07680_),
    .A2(_07686_),
    .B1(_07685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07690_));
 sky130_fd_sc_hd__o211ai_2 _16820_ (.A1(_07684_),
    .A2(_07687_),
    .B1(_07664_),
    .C1(_07665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07691_));
 sky130_fd_sc_hd__o2bb2ai_2 _16821_ (.A1_N(_07664_),
    .A2_N(_07665_),
    .B1(_07688_),
    .B2(_07689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07692_));
 sky130_fd_sc_hd__o2bb2ai_2 _16822_ (.A1_N(_07664_),
    .A2_N(_07665_),
    .B1(_07684_),
    .B2(_07687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07693_));
 sky130_fd_sc_hd__o2111ai_2 _16823_ (.A1(_07680_),
    .A2(_07686_),
    .B1(_07685_),
    .C1(_07664_),
    .D1(_07665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07694_));
 sky130_fd_sc_hd__a21oi_2 _16824_ (.A1(_07693_),
    .A2(_07694_),
    .B1(_07629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07695_));
 sky130_fd_sc_hd__o211ai_2 _16825_ (.A1(_07545_),
    .A2(_07548_),
    .B1(_07691_),
    .C1(_07692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07696_));
 sky130_fd_sc_hd__nand3_2 _16826_ (.A(_07693_),
    .B(_07694_),
    .C(_07629_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07697_));
 sky130_fd_sc_hd__nand2_2 _16827_ (.A(_07696_),
    .B(_07697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07698_));
 sky130_fd_sc_hd__o211ai_2 _16828_ (.A1(_07624_),
    .A2(_07625_),
    .B1(_07696_),
    .C1(_07697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07699_));
 sky130_fd_sc_hd__nand2_2 _16829_ (.A(_07698_),
    .B(_07628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07700_));
 sky130_fd_sc_hd__nand3_2 _16830_ (.A(_07628_),
    .B(_07696_),
    .C(_07697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07701_));
 sky130_fd_sc_hd__a21o_2 _16831_ (.A1(_07696_),
    .A2(_07697_),
    .B1(_07628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07702_));
 sky130_fd_sc_hd__o211ai_2 _16832_ (.A1(_07556_),
    .A2(_07590_),
    .B1(_07699_),
    .C1(_07700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07703_));
 sky130_fd_sc_hd__nand3_2 _16833_ (.A(_07702_),
    .B(_07591_),
    .C(_07701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07704_));
 sky130_fd_sc_hd__nand2_2 _16834_ (.A(_07703_),
    .B(_07704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07705_));
 sky130_fd_sc_hd__nand2_2 _16835_ (.A(\a_l[1] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07706_));
 sky130_fd_sc_hd__a22o_2 _16836_ (.A1(_07473_),
    .A2(_07474_),
    .B1(_07483_),
    .B2(_07487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07707_));
 sky130_fd_sc_hd__and4_2 _16837_ (.A(_07473_),
    .B(_07474_),
    .C(_07483_),
    .D(_07487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07708_));
 sky130_fd_sc_hd__nand4_2 _16838_ (.A(_07473_),
    .B(_07474_),
    .C(_07483_),
    .D(_07487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07709_));
 sky130_fd_sc_hd__a22oi_2 _16839_ (.A1(\a_l[1] ),
    .A2(\b_h[15] ),
    .B1(_07707_),
    .B2(_07709_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07710_));
 sky130_fd_sc_hd__and4_2 _16840_ (.A(_07707_),
    .B(_07709_),
    .C(\a_l[1] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07711_));
 sky130_fd_sc_hd__nor2_2 _16841_ (.A(_07710_),
    .B(_07711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07712_));
 sky130_fd_sc_hd__o211ai_2 _16842_ (.A1(_07710_),
    .A2(_07711_),
    .B1(_07703_),
    .C1(_07704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07713_));
 sky130_fd_sc_hd__nand2_2 _16843_ (.A(_07705_),
    .B(_07712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07714_));
 sky130_fd_sc_hd__o21ai_2 _16844_ (.A1(_07710_),
    .A2(_07711_),
    .B1(_07705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07715_));
 sky130_fd_sc_hd__nand2_2 _16845_ (.A(_07704_),
    .B(_07712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07716_));
 sky130_fd_sc_hd__nand3_2 _16846_ (.A(_07703_),
    .B(_07704_),
    .C(_07712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07717_));
 sky130_fd_sc_hd__nand3_2 _16847_ (.A(_07589_),
    .B(_07713_),
    .C(_07714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07718_));
 sky130_fd_sc_hd__a21oi_2 _16848_ (.A1(_07713_),
    .A2(_07714_),
    .B1(_07589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07719_));
 sky130_fd_sc_hd__nand3_2 _16849_ (.A(_07715_),
    .B(_07717_),
    .C(_07588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07720_));
 sky130_fd_sc_hd__nand2_2 _16850_ (.A(_07718_),
    .B(_07720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07721_));
 sky130_fd_sc_hd__o21ai_2 _16851_ (.A1(_07446_),
    .A2(_07447_),
    .B1(_07444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07722_));
 sky130_fd_sc_hd__inv_2 _16852_ (.A(_07722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07723_));
 sky130_fd_sc_hd__nand2_2 _16853_ (.A(_07721_),
    .B(_07723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07724_));
 sky130_fd_sc_hd__nand3_2 _16854_ (.A(_07718_),
    .B(_07720_),
    .C(_07722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07725_));
 sky130_fd_sc_hd__inv_2 _16855_ (.A(_07725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07726_));
 sky130_fd_sc_hd__o2bb2ai_2 _16856_ (.A1_N(_07424_),
    .A2_N(_07574_),
    .B1(_07569_),
    .B2(_07572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07727_));
 sky130_fd_sc_hd__a21o_2 _16857_ (.A1(_07724_),
    .A2(_07725_),
    .B1(_07727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07728_));
 sky130_fd_sc_hd__nand2_2 _16858_ (.A(_07724_),
    .B(_07727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07729_));
 sky130_fd_sc_hd__nand3_2 _16859_ (.A(_07724_),
    .B(_07727_),
    .C(_07725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07730_));
 sky130_fd_sc_hd__o21a_2 _16860_ (.A1(_07726_),
    .A2(_07729_),
    .B1(_07728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07731_));
 sky130_fd_sc_hd__a31o_2 _16861_ (.A1(_07584_),
    .A2(_07586_),
    .A3(_07731_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07732_));
 sky130_fd_sc_hd__o21ba_2 _16862_ (.A1(_07587_),
    .A2(_07731_),
    .B1_N(_07732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00354_));
 sky130_fd_sc_hd__a32oi_2 _16863_ (.A1(_07693_),
    .A2(_07694_),
    .A3(_07629_),
    .B1(_07627_),
    .B2(_07626_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07733_));
 sky130_fd_sc_hd__o21ai_2 _16864_ (.A1(_07624_),
    .A2(_07625_),
    .B1(_07696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07734_));
 sky130_fd_sc_hd__o21ai_2 _16865_ (.A1(_07628_),
    .A2(_07695_),
    .B1(_07697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07735_));
 sky130_fd_sc_hd__o2bb2ai_2 _16866_ (.A1_N(_07678_),
    .A2_N(_07683_),
    .B1(_07679_),
    .B2(_07674_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07736_));
 sky130_fd_sc_hd__a21oi_2 _16867_ (.A1(_07678_),
    .A2(_07683_),
    .B1(_07680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07737_));
 sky130_fd_sc_hd__nand2_2 _16868_ (.A(\a_l[4] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_2 _16869_ (.A(\a_l[5] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07739_));
 sky130_fd_sc_hd__nand4_2 _16870_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07740_));
 sky130_fd_sc_hd__nand2_2 _16871_ (.A(_07738_),
    .B(_07739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07741_));
 sky130_fd_sc_hd__and4_2 _16872_ (.A(_07741_),
    .B(\b_h[14] ),
    .C(\a_l[3] ),
    .D(_07740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07742_));
 sky130_fd_sc_hd__o2111ai_2 _16873_ (.A1(_02589_),
    .A2(_06605_),
    .B1(\a_l[3] ),
    .C1(\b_h[14] ),
    .D1(_07741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07743_));
 sky130_fd_sc_hd__o2bb2a_2 _16874_ (.A1_N(_07740_),
    .A2_N(_07741_),
    .B1(_09188_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07744_));
 sky130_fd_sc_hd__a22o_2 _16875_ (.A1(\a_l[3] ),
    .A2(\b_h[14] ),
    .B1(_07740_),
    .B2(_07741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07745_));
 sky130_fd_sc_hd__nor2_2 _16876_ (.A(_07742_),
    .B(_07744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07746_));
 sky130_fd_sc_hd__a21o_2 _16877_ (.A1(_07603_),
    .A2(_07606_),
    .B1(_07607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07747_));
 sky130_fd_sc_hd__a21oi_2 _16878_ (.A1(_07603_),
    .A2(_07606_),
    .B1(_07607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07748_));
 sky130_fd_sc_hd__nand2_2 _16879_ (.A(\a_l[6] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07749_));
 sky130_fd_sc_hd__nand2_2 _16880_ (.A(\a_l[7] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07750_));
 sky130_fd_sc_hd__nand2_2 _16881_ (.A(\a_l[8] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07751_));
 sky130_fd_sc_hd__a22oi_2 _16882_ (.A1(\a_l[8] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07752_));
 sky130_fd_sc_hd__nand2_2 _16883_ (.A(_07750_),
    .B(_07751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07753_));
 sky130_fd_sc_hd__nand2_2 _16884_ (.A(\a_l[8] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07754_));
 sky130_fd_sc_hd__nand4_2 _16885_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07755_));
 sky130_fd_sc_hd__o21ai_2 _16886_ (.A1(_02338_),
    .A2(_06867_),
    .B1(_07749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07756_));
 sky130_fd_sc_hd__a21o_2 _16887_ (.A1(_07753_),
    .A2(_07755_),
    .B1(_07749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07757_));
 sky130_fd_sc_hd__o2bb2ai_2 _16888_ (.A1_N(_07753_),
    .A2_N(_07755_),
    .B1(_09231_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07758_));
 sky130_fd_sc_hd__nand3_2 _16889_ (.A(_07755_),
    .B(\b_h[11] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07759_));
 sky130_fd_sc_hd__o211ai_2 _16890_ (.A1(_07752_),
    .A2(_07756_),
    .B1(_07747_),
    .C1(_07757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07760_));
 sky130_fd_sc_hd__o211a_2 _16891_ (.A1(_07759_),
    .A2(_07752_),
    .B1(_07748_),
    .C1(_07758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07761_));
 sky130_fd_sc_hd__o211ai_2 _16892_ (.A1(_07759_),
    .A2(_07752_),
    .B1(_07748_),
    .C1(_07758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07762_));
 sky130_fd_sc_hd__nand2_2 _16893_ (.A(_07760_),
    .B(_07762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07763_));
 sky130_fd_sc_hd__o211ai_2 _16894_ (.A1(_07742_),
    .A2(_07744_),
    .B1(_07760_),
    .C1(_07762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07764_));
 sky130_fd_sc_hd__nand2_2 _16895_ (.A(_07763_),
    .B(_07746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07765_));
 sky130_fd_sc_hd__nand3_2 _16896_ (.A(_07737_),
    .B(_07764_),
    .C(_07765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07766_));
 sky130_fd_sc_hd__a22o_2 _16897_ (.A1(_07743_),
    .A2(_07745_),
    .B1(_07760_),
    .B2(_07762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07767_));
 sky130_fd_sc_hd__and3_2 _16898_ (.A(_07743_),
    .B(_07745_),
    .C(_07760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07768_));
 sky130_fd_sc_hd__nand4_2 _16899_ (.A(_07743_),
    .B(_07745_),
    .C(_07760_),
    .D(_07762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07769_));
 sky130_fd_sc_hd__nand3_2 _16900_ (.A(_07767_),
    .B(_07769_),
    .C(_07736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07770_));
 sky130_fd_sc_hd__nand2_2 _16901_ (.A(_07766_),
    .B(_07770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07771_));
 sky130_fd_sc_hd__a32o_2 _16902_ (.A1(_07600_),
    .A2(_07610_),
    .A3(_07611_),
    .B1(_07599_),
    .B2(_07614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07772_));
 sky130_fd_sc_hd__a21o_2 _16903_ (.A1(_07766_),
    .A2(_07770_),
    .B1(_07772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07773_));
 sky130_fd_sc_hd__nand3_2 _16904_ (.A(_07766_),
    .B(_07770_),
    .C(_07772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_2 _16905_ (.A(_07771_),
    .B(_07772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07775_));
 sky130_fd_sc_hd__nand3b_2 _16906_ (.A_N(_07772_),
    .B(_07770_),
    .C(_07766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_2 _16907_ (.A(_07775_),
    .B(_07776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07777_));
 sky130_fd_sc_hd__nand2_2 _16908_ (.A(_07664_),
    .B(_07690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07778_));
 sky130_fd_sc_hd__o21ai_2 _16909_ (.A1(_07631_),
    .A2(_07663_),
    .B1(_07778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_2 _16910_ (.A(\a_l[9] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_2 _16911_ (.A(\a_l[11] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07781_));
 sky130_fd_sc_hd__a22oi_2 _16912_ (.A1(\a_l[11] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07782_));
 sky130_fd_sc_hd__nand2_2 _16913_ (.A(_07671_),
    .B(_07781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07783_));
 sky130_fd_sc_hd__nand2_2 _16914_ (.A(\a_l[11] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07784_));
 sky130_fd_sc_hd__and4_2 _16915_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07785_));
 sky130_fd_sc_hd__nand4_2 _16916_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07786_));
 sky130_fd_sc_hd__o2111ai_2 _16917_ (.A1(_07668_),
    .A2(_07784_),
    .B1(\a_l[9] ),
    .C1(\b_h[8] ),
    .D1(_07783_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07787_));
 sky130_fd_sc_hd__o2bb2ai_2 _16918_ (.A1_N(_07783_),
    .A2_N(_07786_),
    .B1(_09275_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07788_));
 sky130_fd_sc_hd__nand2_2 _16919_ (.A(_07787_),
    .B(_07788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07789_));
 sky130_fd_sc_hd__nand3_2 _16920_ (.A(_07788_),
    .B(_07633_),
    .C(_07787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07790_));
 sky130_fd_sc_hd__o22a_2 _16921_ (.A1(_09275_),
    .A2(_09613_),
    .B1(_07671_),
    .B2(_07781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07791_));
 sky130_fd_sc_hd__nand2_2 _16922_ (.A(_07780_),
    .B(_07786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07792_));
 sky130_fd_sc_hd__a21oi_2 _16923_ (.A1(_07783_),
    .A2(_07786_),
    .B1(_07780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07793_));
 sky130_fd_sc_hd__a21o_2 _16924_ (.A1(_07783_),
    .A2(_07786_),
    .B1(_07780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07794_));
 sky130_fd_sc_hd__o21ai_2 _16925_ (.A1(_07782_),
    .A2(_07792_),
    .B1(_07634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07795_));
 sky130_fd_sc_hd__o211ai_2 _16926_ (.A1(_07792_),
    .A2(_07782_),
    .B1(_07634_),
    .C1(_07794_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07796_));
 sky130_fd_sc_hd__o21ai_2 _16927_ (.A1(_07793_),
    .A2(_07795_),
    .B1(_07790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07797_));
 sky130_fd_sc_hd__o31a_2 _16928_ (.A1(_09253_),
    .A2(_09613_),
    .A3(_07669_),
    .B1(_07672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07798_));
 sky130_fd_sc_hd__a21oi_2 _16929_ (.A1(_07667_),
    .A2(_07672_),
    .B1(_07669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07799_));
 sky130_fd_sc_hd__o211a_2 _16930_ (.A1(_07793_),
    .A2(_07795_),
    .B1(_07798_),
    .C1(_07790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07800_));
 sky130_fd_sc_hd__a21oi_2 _16931_ (.A1(_07790_),
    .A2(_07796_),
    .B1(_07798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07801_));
 sky130_fd_sc_hd__nand2_2 _16932_ (.A(_07797_),
    .B(_07798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07802_));
 sky130_fd_sc_hd__o21ai_2 _16933_ (.A1(_07793_),
    .A2(_07795_),
    .B1(_07799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07803_));
 sky130_fd_sc_hd__o211ai_2 _16934_ (.A1(_07793_),
    .A2(_07795_),
    .B1(_07799_),
    .C1(_07790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07804_));
 sky130_fd_sc_hd__nand2_2 _16935_ (.A(_07802_),
    .B(_07804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07805_));
 sky130_fd_sc_hd__a31o_2 _16936_ (.A1(_07649_),
    .A2(_07650_),
    .A3(_07637_),
    .B1(_07636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07806_));
 sky130_fd_sc_hd__a21boi_2 _16937_ (.A1(_07656_),
    .A2(_07636_),
    .B1_N(_07655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07807_));
 sky130_fd_sc_hd__a21o_2 _16938_ (.A1(_07641_),
    .A2(_07642_),
    .B1(_07640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07808_));
 sky130_fd_sc_hd__nand2_2 _16939_ (.A(\a_l[15] ),
    .B(\b_h[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07809_));
 sky130_fd_sc_hd__nand2_2 _16940_ (.A(_07645_),
    .B(_07809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07810_));
 sky130_fd_sc_hd__nand2_2 _16941_ (.A(\a_l[15] ),
    .B(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07811_));
 sky130_fd_sc_hd__nand4_2 _16942_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[2] ),
    .D(\b_h[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_2 _16943_ (.A(_07810_),
    .B(_07812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07813_));
 sky130_fd_sc_hd__o21ai_2 _16944_ (.A1(_07640_),
    .A2(_07643_),
    .B1(_07813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07814_));
 sky130_fd_sc_hd__o211ai_2 _16945_ (.A1(_07640_),
    .A2(_07643_),
    .B1(_07647_),
    .C1(_07813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07815_));
 sky130_fd_sc_hd__nand3_2 _16946_ (.A(_07644_),
    .B(_07810_),
    .C(_07812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07816_));
 sky130_fd_sc_hd__nand4_2 _16947_ (.A(_07644_),
    .B(_07653_),
    .C(_07810_),
    .D(_07812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07817_));
 sky130_fd_sc_hd__nand2_2 _16948_ (.A(_07815_),
    .B(_07817_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07818_));
 sky130_fd_sc_hd__a22oi_2 _16949_ (.A1(\a_l[13] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07819_));
 sky130_fd_sc_hd__a22o_2 _16950_ (.A1(\a_l[13] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07820_));
 sky130_fd_sc_hd__nand2_2 _16951_ (.A(\a_l[13] ),
    .B(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07821_));
 sky130_fd_sc_hd__and4_2 _16952_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07822_));
 sky130_fd_sc_hd__nor2_2 _16953_ (.A(_07819_),
    .B(_07822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07823_));
 sky130_fd_sc_hd__o21ai_2 _16954_ (.A1(_07113_),
    .A2(_07821_),
    .B1(_07820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07824_));
 sky130_fd_sc_hd__o21ai_2 _16955_ (.A1(_07819_),
    .A2(_07822_),
    .B1(_07818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07825_));
 sky130_fd_sc_hd__o211ai_2 _16956_ (.A1(_07652_),
    .A2(_07816_),
    .B1(_07823_),
    .C1(_07815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07826_));
 sky130_fd_sc_hd__nand2_2 _16957_ (.A(_07818_),
    .B(_07823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07827_));
 sky130_fd_sc_hd__o211ai_2 _16958_ (.A1(_07652_),
    .A2(_07816_),
    .B1(_07824_),
    .C1(_07815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_2 _16959_ (.A(_07825_),
    .B(_07826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07829_));
 sky130_fd_sc_hd__nand4_2 _16960_ (.A(_07656_),
    .B(_07806_),
    .C(_07825_),
    .D(_07826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07830_));
 sky130_fd_sc_hd__nand4_2 _16961_ (.A(_07655_),
    .B(_07658_),
    .C(_07827_),
    .D(_07828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07831_));
 sky130_fd_sc_hd__nand2_2 _16962_ (.A(_07830_),
    .B(_07831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07832_));
 sky130_fd_sc_hd__o21ai_2 _16963_ (.A1(_07800_),
    .A2(_07801_),
    .B1(_07831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07833_));
 sky130_fd_sc_hd__o211a_2 _16964_ (.A1(_07800_),
    .A2(_07801_),
    .B1(_07830_),
    .C1(_07831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07834_));
 sky130_fd_sc_hd__o211ai_2 _16965_ (.A1(_07800_),
    .A2(_07801_),
    .B1(_07830_),
    .C1(_07831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07835_));
 sky130_fd_sc_hd__nand2_2 _16966_ (.A(_07832_),
    .B(_07805_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07836_));
 sky130_fd_sc_hd__o2bb2ai_2 _16967_ (.A1_N(_07802_),
    .A2_N(_07804_),
    .B1(_07807_),
    .B2(_07829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07837_));
 sky130_fd_sc_hd__nand3_2 _16968_ (.A(_07805_),
    .B(_07830_),
    .C(_07831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07838_));
 sky130_fd_sc_hd__o21ai_2 _16969_ (.A1(_07800_),
    .A2(_07801_),
    .B1(_07832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07839_));
 sky130_fd_sc_hd__nand2_2 _16970_ (.A(_07835_),
    .B(_07836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07840_));
 sky130_fd_sc_hd__o211ai_2 _16971_ (.A1(_07631_),
    .A2(_07663_),
    .B1(_07778_),
    .C1(_07836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07841_));
 sky130_fd_sc_hd__nand4_2 _16972_ (.A(_07665_),
    .B(_07778_),
    .C(_07835_),
    .D(_07836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07842_));
 sky130_fd_sc_hd__nand3_2 _16973_ (.A(_07779_),
    .B(_07838_),
    .C(_07839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07843_));
 sky130_fd_sc_hd__a22oi_2 _16974_ (.A1(_07775_),
    .A2(_07776_),
    .B1(_07840_),
    .B2(_07779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07844_));
 sky130_fd_sc_hd__o211a_2 _16975_ (.A1(_07834_),
    .A2(_07841_),
    .B1(_07843_),
    .C1(_07777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07845_));
 sky130_fd_sc_hd__o211ai_2 _16976_ (.A1(_07834_),
    .A2(_07841_),
    .B1(_07843_),
    .C1(_07777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07846_));
 sky130_fd_sc_hd__a22oi_2 _16977_ (.A1(_07773_),
    .A2(_07774_),
    .B1(_07842_),
    .B2(_07843_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07847_));
 sky130_fd_sc_hd__a21o_2 _16978_ (.A1(_07842_),
    .A2(_07843_),
    .B1(_07777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07848_));
 sky130_fd_sc_hd__a221oi_2 _16979_ (.A1(_07844_),
    .A2(_07842_),
    .B1(_07734_),
    .B2(_07697_),
    .C1(_07847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07849_));
 sky130_fd_sc_hd__nand3_2 _16980_ (.A(_07735_),
    .B(_07846_),
    .C(_07848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07850_));
 sky130_fd_sc_hd__a2bb2oi_2 _16981_ (.A1_N(_07695_),
    .A2_N(_07733_),
    .B1(_07846_),
    .B2(_07848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07851_));
 sky130_fd_sc_hd__o22ai_2 _16982_ (.A1(_07695_),
    .A2(_07733_),
    .B1(_07845_),
    .B2(_07847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07852_));
 sky130_fd_sc_hd__a31o_2 _16983_ (.A1(_07593_),
    .A2(\b_h[14] ),
    .A3(\a_l[2] ),
    .B1(_07594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07853_));
 sky130_fd_sc_hd__nand2_2 _16984_ (.A(_07620_),
    .B(_07622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07854_));
 sky130_fd_sc_hd__and3_2 _16985_ (.A(_07621_),
    .B(_07853_),
    .C(_07854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07855_));
 sky130_fd_sc_hd__nand3_2 _16986_ (.A(_07621_),
    .B(_07853_),
    .C(_07854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07856_));
 sky130_fd_sc_hd__a21o_2 _16987_ (.A1(_07621_),
    .A2(_07854_),
    .B1(_07853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07857_));
 sky130_fd_sc_hd__nand4_2 _16988_ (.A(_07857_),
    .B(\b_h[15] ),
    .C(\a_l[2] ),
    .D(_07856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07858_));
 sky130_fd_sc_hd__a22o_2 _16989_ (.A1(\a_l[2] ),
    .A2(\b_h[15] ),
    .B1(_07856_),
    .B2(_07857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07859_));
 sky130_fd_sc_hd__nand2_2 _16990_ (.A(_07858_),
    .B(_07859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07860_));
 sky130_fd_sc_hd__nand3_2 _16991_ (.A(_07850_),
    .B(_07852_),
    .C(_07860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07861_));
 sky130_fd_sc_hd__o21bai_2 _16992_ (.A1(_07849_),
    .A2(_07851_),
    .B1_N(_07860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07862_));
 sky130_fd_sc_hd__o21ai_2 _16993_ (.A1(_07849_),
    .A2(_07851_),
    .B1(_07860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07863_));
 sky130_fd_sc_hd__nand4_2 _16994_ (.A(_07850_),
    .B(_07852_),
    .C(_07858_),
    .D(_07859_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07864_));
 sky130_fd_sc_hd__nand2_2 _16995_ (.A(_07703_),
    .B(_07716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07865_));
 sky130_fd_sc_hd__a21boi_2 _16996_ (.A1(_07704_),
    .A2(_07712_),
    .B1_N(_07703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07866_));
 sky130_fd_sc_hd__a21oi_2 _16997_ (.A1(_07863_),
    .A2(_07864_),
    .B1(_07865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07867_));
 sky130_fd_sc_hd__nand3_2 _16998_ (.A(_07861_),
    .B(_07862_),
    .C(_07866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07868_));
 sky130_fd_sc_hd__nand3_2 _16999_ (.A(_07863_),
    .B(_07865_),
    .C(_07864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07869_));
 sky130_fd_sc_hd__o21ai_2 _17000_ (.A1(_07706_),
    .A2(_07708_),
    .B1(_07707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07870_));
 sky130_fd_sc_hd__o21a_2 _17001_ (.A1(_07706_),
    .A2(_07708_),
    .B1(_07707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07871_));
 sky130_fd_sc_hd__a21o_2 _17002_ (.A1(_07868_),
    .A2(_07869_),
    .B1(_07871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07872_));
 sky130_fd_sc_hd__o2111ai_2 _17003_ (.A1(_07708_),
    .A2(_07706_),
    .B1(_07707_),
    .C1(_07868_),
    .D1(_07869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07873_));
 sky130_fd_sc_hd__a21oi_2 _17004_ (.A1(_07868_),
    .A2(_07869_),
    .B1(_07870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07874_));
 sky130_fd_sc_hd__a21o_2 _17005_ (.A1(_07868_),
    .A2(_07869_),
    .B1(_07870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07875_));
 sky130_fd_sc_hd__nand3_2 _17006_ (.A(_07868_),
    .B(_07869_),
    .C(_07870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07876_));
 sky130_fd_sc_hd__a31oi_2 _17007_ (.A1(_07589_),
    .A2(_07713_),
    .A3(_07714_),
    .B1(_07723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07877_));
 sky130_fd_sc_hd__o21ai_2 _17008_ (.A1(_07722_),
    .A2(_07719_),
    .B1(_07718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07878_));
 sky130_fd_sc_hd__nand3_2 _17009_ (.A(_07872_),
    .B(_07878_),
    .C(_07873_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07879_));
 sky130_fd_sc_hd__o211ai_2 _17010_ (.A1(_07722_),
    .A2(_07719_),
    .B1(_07718_),
    .C1(_07876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07880_));
 sky130_fd_sc_hd__o211ai_2 _17011_ (.A1(_07719_),
    .A2(_07877_),
    .B1(_07876_),
    .C1(_07875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07881_));
 sky130_fd_sc_hd__o21ai_2 _17012_ (.A1(_07874_),
    .A2(_07880_),
    .B1(_07879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07882_));
 sky130_fd_sc_hd__o2bb2a_2 _17013_ (.A1_N(_07587_),
    .A2_N(_07728_),
    .B1(_07729_),
    .B2(_07726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07883_));
 sky130_fd_sc_hd__a21oi_2 _17014_ (.A1(_07882_),
    .A2(_07883_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07884_));
 sky130_fd_sc_hd__o21a_2 _17015_ (.A1(_07882_),
    .A2(_07883_),
    .B1(_07884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00355_));
 sky130_fd_sc_hd__a31oi_2 _17016_ (.A1(_07863_),
    .A2(_07865_),
    .A3(_07864_),
    .B1(_07870_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07885_));
 sky130_fd_sc_hd__nand2_2 _17017_ (.A(_07869_),
    .B(_07871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07886_));
 sky130_fd_sc_hd__nor2_2 _17018_ (.A(_09188_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07887_));
 sky130_fd_sc_hd__a31o_2 _17019_ (.A1(\a_l[4] ),
    .A2(\a_l[5] ),
    .A3(_02588_),
    .B1(_07742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07888_));
 sky130_fd_sc_hd__nand2_2 _17020_ (.A(_07766_),
    .B(_07772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07889_));
 sky130_fd_sc_hd__a22oi_2 _17021_ (.A1(_07740_),
    .A2(_07743_),
    .B1(_07770_),
    .B2(_07889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07890_));
 sky130_fd_sc_hd__and3b_2 _17022_ (.A_N(_07888_),
    .B(_07889_),
    .C(_07770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07891_));
 sky130_fd_sc_hd__o2111ai_2 _17023_ (.A1(_02589_),
    .A2(_06605_),
    .B1(_07743_),
    .C1(_07770_),
    .D1(_07774_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07892_));
 sky130_fd_sc_hd__o22ai_2 _17024_ (.A1(_09188_),
    .A2(_09679_),
    .B1(_07890_),
    .B2(_07891_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07893_));
 sky130_fd_sc_hd__nand3b_2 _17025_ (.A_N(_07890_),
    .B(_07892_),
    .C(_07887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07894_));
 sky130_fd_sc_hd__nand2_2 _17026_ (.A(_07893_),
    .B(_07894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07895_));
 sky130_fd_sc_hd__a2bb2oi_2 _17027_ (.A1_N(_07834_),
    .A2_N(_07841_),
    .B1(_07843_),
    .B2(_07777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07896_));
 sky130_fd_sc_hd__o2bb2ai_2 _17028_ (.A1_N(_07777_),
    .A2_N(_07843_),
    .B1(_07841_),
    .B2(_07834_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07897_));
 sky130_fd_sc_hd__a31oi_2 _17029_ (.A1(_07647_),
    .A2(_07808_),
    .A3(_07813_),
    .B1(_07824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07898_));
 sky130_fd_sc_hd__a21oi_2 _17030_ (.A1(\a_l[14] ),
    .A2(\b_h[2] ),
    .B1(_07811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07899_));
 sky130_fd_sc_hd__nand3_2 _17031_ (.A(_07642_),
    .B(\b_h[3] ),
    .C(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07900_));
 sky130_fd_sc_hd__a22o_2 _17032_ (.A1(\a_l[14] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07901_));
 sky130_fd_sc_hd__and4_2 _17033_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07902_));
 sky130_fd_sc_hd__nand4_2 _17034_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07903_));
 sky130_fd_sc_hd__nand3_2 _17035_ (.A(_07392_),
    .B(\b_h[5] ),
    .C(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07904_));
 sky130_fd_sc_hd__nand3_2 _17036_ (.A(_07821_),
    .B(\b_h[4] ),
    .C(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07905_));
 sky130_fd_sc_hd__nand3_2 _17037_ (.A(_07899_),
    .B(_07901_),
    .C(_07903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07906_));
 sky130_fd_sc_hd__inv_2 _17038_ (.A(_07906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07907_));
 sky130_fd_sc_hd__a21o_2 _17039_ (.A1(_07901_),
    .A2(_07903_),
    .B1(_07899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07908_));
 sky130_fd_sc_hd__nand3_2 _17040_ (.A(_07900_),
    .B(_07901_),
    .C(_07903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07909_));
 sky130_fd_sc_hd__nand3_2 _17041_ (.A(_07899_),
    .B(_07904_),
    .C(_07905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07910_));
 sky130_fd_sc_hd__nand2_2 _17042_ (.A(_07909_),
    .B(_07910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07911_));
 sky130_fd_sc_hd__nand3_2 _17043_ (.A(_07817_),
    .B(_07909_),
    .C(_07910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07912_));
 sky130_fd_sc_hd__o22ai_2 _17044_ (.A1(_07819_),
    .A2(_07822_),
    .B1(_07652_),
    .B2(_07816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07913_));
 sky130_fd_sc_hd__a22oi_2 _17045_ (.A1(_07906_),
    .A2(_07908_),
    .B1(_07913_),
    .B2(_07815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07914_));
 sky130_fd_sc_hd__o211a_2 _17046_ (.A1(_07646_),
    .A2(_07814_),
    .B1(_07911_),
    .C1(_07913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07915_));
 sky130_fd_sc_hd__o211ai_2 _17047_ (.A1(_07646_),
    .A2(_07814_),
    .B1(_07911_),
    .C1(_07913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07916_));
 sky130_fd_sc_hd__o21a_2 _17048_ (.A1(_07898_),
    .A2(_07912_),
    .B1(_07916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07917_));
 sky130_fd_sc_hd__o21ai_2 _17049_ (.A1(_07912_),
    .A2(_07898_),
    .B1(_07916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07918_));
 sky130_fd_sc_hd__and3_2 _17050_ (.A(_07783_),
    .B(\b_h[8] ),
    .C(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07919_));
 sky130_fd_sc_hd__a31o_2 _17051_ (.A1(\a_l[9] ),
    .A2(_07783_),
    .A3(\b_h[8] ),
    .B1(_07785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07920_));
 sky130_fd_sc_hd__and2_2 _17052_ (.A(\a_l[10] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07921_));
 sky130_fd_sc_hd__nand2_2 _17053_ (.A(\a_l[10] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_2 _17054_ (.A(\a_l[12] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07923_));
 sky130_fd_sc_hd__nand2_2 _17055_ (.A(_07784_),
    .B(_07923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07924_));
 sky130_fd_sc_hd__nand2_2 _17056_ (.A(\a_l[12] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07925_));
 sky130_fd_sc_hd__and4_2 _17057_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07926_));
 sky130_fd_sc_hd__nand4_2 _17058_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07927_));
 sky130_fd_sc_hd__and3_2 _17059_ (.A(_07924_),
    .B(_07927_),
    .C(_07921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07928_));
 sky130_fd_sc_hd__o2111ai_2 _17060_ (.A1(_07781_),
    .A2(_07925_),
    .B1(\a_l[10] ),
    .C1(\b_h[8] ),
    .D1(_07924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07929_));
 sky130_fd_sc_hd__a21o_2 _17061_ (.A1(_07924_),
    .A2(_07927_),
    .B1(_07921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07930_));
 sky130_fd_sc_hd__o221ai_2 _17062_ (.A1(_09286_),
    .A2(_09613_),
    .B1(_07781_),
    .B2(_07925_),
    .C1(_07924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07931_));
 sky130_fd_sc_hd__a21o_2 _17063_ (.A1(_07924_),
    .A2(_07927_),
    .B1(_07922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07932_));
 sky130_fd_sc_hd__nand2_2 _17064_ (.A(_07930_),
    .B(_07822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07933_));
 sky130_fd_sc_hd__nand3_2 _17065_ (.A(_07930_),
    .B(_07822_),
    .C(_07929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07934_));
 sky130_fd_sc_hd__o211ai_2 _17066_ (.A1(_07244_),
    .A2(_07632_),
    .B1(_07931_),
    .C1(_07932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07935_));
 sky130_fd_sc_hd__a2bb2oi_2 _17067_ (.A1_N(_07782_),
    .A2_N(_07791_),
    .B1(_07934_),
    .B2(_07935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07936_));
 sky130_fd_sc_hd__a22o_2 _17068_ (.A1(_07783_),
    .A2(_07792_),
    .B1(_07934_),
    .B2(_07935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07937_));
 sky130_fd_sc_hd__o211a_2 _17069_ (.A1(_07785_),
    .A2(_07919_),
    .B1(_07934_),
    .C1(_07935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07938_));
 sky130_fd_sc_hd__o211ai_2 _17070_ (.A1(_07785_),
    .A2(_07919_),
    .B1(_07934_),
    .C1(_07935_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07939_));
 sky130_fd_sc_hd__o22ai_2 _17071_ (.A1(_07914_),
    .A2(_07915_),
    .B1(_07936_),
    .B2(_07938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07940_));
 sky130_fd_sc_hd__o21ai_2 _17072_ (.A1(_07898_),
    .A2(_07912_),
    .B1(_07939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07941_));
 sky130_fd_sc_hd__o211ai_2 _17073_ (.A1(_07898_),
    .A2(_07912_),
    .B1(_07916_),
    .C1(_07939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07942_));
 sky130_fd_sc_hd__nand3_2 _17074_ (.A(_07917_),
    .B(_07937_),
    .C(_07939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07943_));
 sky130_fd_sc_hd__o21ai_2 _17075_ (.A1(_07936_),
    .A2(_07938_),
    .B1(_07917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07944_));
 sky130_fd_sc_hd__nand3_2 _17076_ (.A(_07918_),
    .B(_07937_),
    .C(_07939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07945_));
 sky130_fd_sc_hd__o21ai_2 _17077_ (.A1(_07936_),
    .A2(_07942_),
    .B1(_07940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07946_));
 sky130_fd_sc_hd__nand4_2 _17078_ (.A(_07830_),
    .B(_07833_),
    .C(_07944_),
    .D(_07945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07947_));
 sky130_fd_sc_hd__o21ai_2 _17079_ (.A1(_07634_),
    .A2(_07789_),
    .B1(_07803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07948_));
 sky130_fd_sc_hd__o21ai_2 _17080_ (.A1(_07749_),
    .A2(_07752_),
    .B1(_07755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07949_));
 sky130_fd_sc_hd__o22a_2 _17081_ (.A1(_02338_),
    .A2(_06867_),
    .B1(_07749_),
    .B2(_07752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07950_));
 sky130_fd_sc_hd__and2_2 _17082_ (.A(\a_l[7] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07951_));
 sky130_fd_sc_hd__nand2_2 _17083_ (.A(\a_l[7] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07952_));
 sky130_fd_sc_hd__nand2_2 _17084_ (.A(\a_l[9] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07953_));
 sky130_fd_sc_hd__nand2_2 _17085_ (.A(_07754_),
    .B(_07953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07954_));
 sky130_fd_sc_hd__nand4_2 _17086_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07955_));
 sky130_fd_sc_hd__o221ai_2 _17087_ (.A1(_09242_),
    .A2(_09646_),
    .B1(_02338_),
    .B2(_06985_),
    .C1(_07954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07956_));
 sky130_fd_sc_hd__a21o_2 _17088_ (.A1(_07954_),
    .A2(_07955_),
    .B1(_07952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07957_));
 sky130_fd_sc_hd__o2bb2a_2 _17089_ (.A1_N(_07954_),
    .A2_N(_07955_),
    .B1(_09242_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07958_));
 sky130_fd_sc_hd__a22o_2 _17090_ (.A1(\a_l[7] ),
    .A2(\b_h[11] ),
    .B1(_07954_),
    .B2(_07955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07959_));
 sky130_fd_sc_hd__o311a_2 _17091_ (.A1(_09253_),
    .A2(_09275_),
    .A3(_02338_),
    .B1(_07951_),
    .C1(_07954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07960_));
 sky130_fd_sc_hd__o2111ai_2 _17092_ (.A1(_02338_),
    .A2(_06985_),
    .B1(\a_l[7] ),
    .C1(\b_h[11] ),
    .D1(_07954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07961_));
 sky130_fd_sc_hd__o221a_2 _17093_ (.A1(_07749_),
    .A2(_07752_),
    .B1(_07958_),
    .B2(_07960_),
    .C1(_07755_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07962_));
 sky130_fd_sc_hd__nand3_2 _17094_ (.A(_07950_),
    .B(_07956_),
    .C(_07957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07963_));
 sky130_fd_sc_hd__nand3_2 _17095_ (.A(_07959_),
    .B(_07961_),
    .C(_07949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07964_));
 sky130_fd_sc_hd__inv_2 _17096_ (.A(_07964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_2 _17097_ (.A(\a_l[4] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07966_));
 sky130_fd_sc_hd__a22oi_2 _17098_ (.A1(\a_l[6] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07967_));
 sky130_fd_sc_hd__and4_2 _17099_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07968_));
 sky130_fd_sc_hd__a21oi_2 _17100_ (.A1(\a_l[4] ),
    .A2(\b_h[14] ),
    .B1(_07968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07969_));
 sky130_fd_sc_hd__a41o_2 _17101_ (.A1(\a_l[5] ),
    .A2(\a_l[6] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_07966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07970_));
 sky130_fd_sc_hd__nor2_2 _17102_ (.A(_07967_),
    .B(_07970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07971_));
 sky130_fd_sc_hd__o22a_2 _17103_ (.A1(_09199_),
    .A2(_09668_),
    .B1(_07967_),
    .B2(_07968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07972_));
 sky130_fd_sc_hd__o21ai_2 _17104_ (.A1(_07967_),
    .A2(_07968_),
    .B1(_07966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07973_));
 sky130_fd_sc_hd__o21ai_2 _17105_ (.A1(_07967_),
    .A2(_07970_),
    .B1(_07973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07974_));
 sky130_fd_sc_hd__o21a_2 _17106_ (.A1(_07967_),
    .A2(_07970_),
    .B1(_07973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07975_));
 sky130_fd_sc_hd__o2bb2ai_2 _17107_ (.A1_N(_07963_),
    .A2_N(_07964_),
    .B1(_07971_),
    .B2(_07972_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07976_));
 sky130_fd_sc_hd__o2111ai_2 _17108_ (.A1(_07967_),
    .A2(_07970_),
    .B1(_07973_),
    .C1(_07964_),
    .D1(_07963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07977_));
 sky130_fd_sc_hd__nand3_2 _17109_ (.A(_07976_),
    .B(_07977_),
    .C(_07948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07978_));
 sky130_fd_sc_hd__nand3_2 _17110_ (.A(_07963_),
    .B(_07964_),
    .C(_07974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07979_));
 sky130_fd_sc_hd__a21oi_2 _17111_ (.A1(_07963_),
    .A2(_07964_),
    .B1(_07974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07980_));
 sky130_fd_sc_hd__o211ai_2 _17112_ (.A1(_07634_),
    .A2(_07789_),
    .B1(_07803_),
    .C1(_07979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07981_));
 sky130_fd_sc_hd__a21o_2 _17113_ (.A1(_07976_),
    .A2(_07977_),
    .B1(_07948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_07982_));
 sky130_fd_sc_hd__o21ai_2 _17114_ (.A1(_07980_),
    .A2(_07981_),
    .B1(_07978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07983_));
 sky130_fd_sc_hd__o21ai_2 _17115_ (.A1(_07746_),
    .A2(_07761_),
    .B1(_07760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07984_));
 sky130_fd_sc_hd__o22ai_2 _17116_ (.A1(_07761_),
    .A2(_07768_),
    .B1(_07980_),
    .B2(_07981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07985_));
 sky130_fd_sc_hd__o211ai_2 _17117_ (.A1(_07761_),
    .A2(_07768_),
    .B1(_07978_),
    .C1(_07982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07986_));
 sky130_fd_sc_hd__nand2_2 _17118_ (.A(_07983_),
    .B(_07984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07987_));
 sky130_fd_sc_hd__nand2_2 _17119_ (.A(_07986_),
    .B(_07987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07988_));
 sky130_fd_sc_hd__a21oi_2 _17120_ (.A1(_07830_),
    .A2(_07833_),
    .B1(_07946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07989_));
 sky130_fd_sc_hd__nand4_2 _17121_ (.A(_07831_),
    .B(_07837_),
    .C(_07940_),
    .D(_07943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07990_));
 sky130_fd_sc_hd__o211ai_2 _17122_ (.A1(_07983_),
    .A2(_07984_),
    .B1(_07987_),
    .C1(_07947_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07991_));
 sky130_fd_sc_hd__nand2_2 _17123_ (.A(_07990_),
    .B(_07991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07992_));
 sky130_fd_sc_hd__a31oi_2 _17124_ (.A1(_07947_),
    .A2(_07986_),
    .A3(_07987_),
    .B1(_07989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07993_));
 sky130_fd_sc_hd__nand2_2 _17125_ (.A(_07947_),
    .B(_07990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07994_));
 sky130_fd_sc_hd__nand4_2 _17126_ (.A(_07947_),
    .B(_07986_),
    .C(_07987_),
    .D(_07990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07995_));
 sky130_fd_sc_hd__nand2_2 _17127_ (.A(_07994_),
    .B(_07988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07996_));
 sky130_fd_sc_hd__o21ai_2 _17128_ (.A1(_07989_),
    .A2(_07991_),
    .B1(_07996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07997_));
 sky130_fd_sc_hd__nor2_2 _17129_ (.A(_07896_),
    .B(_07997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07998_));
 sky130_fd_sc_hd__o211ai_2 _17130_ (.A1(_07989_),
    .A2(_07991_),
    .B1(_07996_),
    .C1(_07897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_07999_));
 sky130_fd_sc_hd__a21oi_2 _17131_ (.A1(_07995_),
    .A2(_07996_),
    .B1(_07897_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08000_));
 sky130_fd_sc_hd__o21bai_2 _17132_ (.A1(_07998_),
    .A2(_08000_),
    .B1_N(_07895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08001_));
 sky130_fd_sc_hd__nand3b_2 _17133_ (.A_N(_08000_),
    .B(_07895_),
    .C(_07999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08002_));
 sky130_fd_sc_hd__a21oi_2 _17134_ (.A1(_07896_),
    .A2(_07997_),
    .B1(_07895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08003_));
 sky130_fd_sc_hd__o21ai_2 _17135_ (.A1(_07896_),
    .A2(_07997_),
    .B1(_08003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08004_));
 sky130_fd_sc_hd__o21ai_2 _17136_ (.A1(_07998_),
    .A2(_08000_),
    .B1(_07895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08005_));
 sky130_fd_sc_hd__a21o_2 _17137_ (.A1(_07850_),
    .A2(_07860_),
    .B1(_07851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08006_));
 sky130_fd_sc_hd__a21oi_2 _17138_ (.A1(_07850_),
    .A2(_07860_),
    .B1(_07851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08007_));
 sky130_fd_sc_hd__a21oi_2 _17139_ (.A1(_08004_),
    .A2(_08005_),
    .B1(_08007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08008_));
 sky130_fd_sc_hd__nand3_2 _17140_ (.A(_08006_),
    .B(_08002_),
    .C(_08001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08009_));
 sky130_fd_sc_hd__a21oi_2 _17141_ (.A1(_08001_),
    .A2(_08002_),
    .B1(_08006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08010_));
 sky130_fd_sc_hd__nand3_2 _17142_ (.A(_08004_),
    .B(_08005_),
    .C(_08007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_2 _17143_ (.A(_08009_),
    .B(_08011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08012_));
 sky130_fd_sc_hd__a31o_2 _17144_ (.A1(_07857_),
    .A2(\b_h[15] ),
    .A3(\a_l[2] ),
    .B1(_07855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08013_));
 sky130_fd_sc_hd__a31oi_2 _17145_ (.A1(_07857_),
    .A2(\b_h[15] ),
    .A3(\a_l[2] ),
    .B1(_07855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08014_));
 sky130_fd_sc_hd__nand3_2 _17146_ (.A(_08009_),
    .B(_08011_),
    .C(_08014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08015_));
 sky130_fd_sc_hd__nand2_2 _17147_ (.A(_08012_),
    .B(_08013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08016_));
 sky130_fd_sc_hd__a21oi_2 _17148_ (.A1(_08009_),
    .A2(_08011_),
    .B1(_08013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08017_));
 sky130_fd_sc_hd__nand3_2 _17149_ (.A(_08009_),
    .B(_08011_),
    .C(_08013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08018_));
 sky130_fd_sc_hd__nand3_2 _17150_ (.A(_07868_),
    .B(_07886_),
    .C(_08018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08019_));
 sky130_fd_sc_hd__a21o_2 _17151_ (.A1(_08012_),
    .A2(_08014_),
    .B1(_08019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08020_));
 sky130_fd_sc_hd__o211ai_2 _17152_ (.A1(_07867_),
    .A2(_07885_),
    .B1(_08015_),
    .C1(_08016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08021_));
 sky130_fd_sc_hd__o21a_2 _17153_ (.A1(_08017_),
    .A2(_08019_),
    .B1(_08021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08022_));
 sky130_fd_sc_hd__o21ai_2 _17154_ (.A1(_08017_),
    .A2(_08019_),
    .B1(_08021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08023_));
 sky130_fd_sc_hd__o2111a_2 _17155_ (.A1(_07726_),
    .A2(_07729_),
    .B1(_07879_),
    .C1(_07881_),
    .D1(_07728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08024_));
 sky130_fd_sc_hd__nand4_2 _17156_ (.A(_07728_),
    .B(_07730_),
    .C(_07879_),
    .D(_07881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08025_));
 sky130_fd_sc_hd__o21ai_2 _17157_ (.A1(_07874_),
    .A2(_07880_),
    .B1(_07730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08026_));
 sky130_fd_sc_hd__a21boi_2 _17158_ (.A1(_07730_),
    .A2(_07881_),
    .B1_N(_07879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08027_));
 sky130_fd_sc_hd__a31o_2 _17159_ (.A1(_07584_),
    .A2(_07586_),
    .A3(_08024_),
    .B1(_08027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08028_));
 sky130_fd_sc_hd__a311o_2 _17160_ (.A1(_07584_),
    .A2(_08024_),
    .A3(_07586_),
    .B1(_08022_),
    .C1(_08027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08029_));
 sky130_fd_sc_hd__nand2_2 _17161_ (.A(_08028_),
    .B(_08022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08030_));
 sky130_fd_sc_hd__and3_2 _17162_ (.A(_09690_),
    .B(_08029_),
    .C(_08030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00356_));
 sky130_fd_sc_hd__o2bb2a_2 _17163_ (.A1_N(_07893_),
    .A2_N(_07894_),
    .B1(_07896_),
    .B2(_07997_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08031_));
 sky130_fd_sc_hd__nand2_2 _17164_ (.A(\a_l[4] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08032_));
 sky130_fd_sc_hd__nor2_2 _17165_ (.A(_07967_),
    .B(_07969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08033_));
 sky130_fd_sc_hd__nand2_2 _17166_ (.A(_07978_),
    .B(_07984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08034_));
 sky130_fd_sc_hd__o211ai_2 _17167_ (.A1(_07980_),
    .A2(_07981_),
    .B1(_08033_),
    .C1(_08034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08035_));
 sky130_fd_sc_hd__o211ai_2 _17168_ (.A1(_07967_),
    .A2(_07969_),
    .B1(_07978_),
    .C1(_07985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08036_));
 sky130_fd_sc_hd__a21o_2 _17169_ (.A1(_08035_),
    .A2(_08036_),
    .B1(_08032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08037_));
 sky130_fd_sc_hd__a32o_2 _17170_ (.A1(_07982_),
    .A2(_08034_),
    .A3(_08033_),
    .B1(\a_l[4] ),
    .B2(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08038_));
 sky130_fd_sc_hd__o211ai_2 _17171_ (.A1(_09199_),
    .A2(_09679_),
    .B1(_08035_),
    .C1(_08036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08039_));
 sky130_fd_sc_hd__nand2_2 _17172_ (.A(_08037_),
    .B(_08039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08040_));
 sky130_fd_sc_hd__nor2_2 _17173_ (.A(_09373_),
    .B(_09602_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08041_));
 sky130_fd_sc_hd__and4_2 _17174_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08042_));
 sky130_fd_sc_hd__nand4_2 _17175_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[4] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08043_));
 sky130_fd_sc_hd__a22o_2 _17176_ (.A1(\a_l[15] ),
    .A2(\b_h[4] ),
    .B1(\b_h[5] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08044_));
 sky130_fd_sc_hd__nand2_2 _17177_ (.A(_08043_),
    .B(_08044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08045_));
 sky130_fd_sc_hd__o31a_2 _17178_ (.A1(_09373_),
    .A2(_09592_),
    .A3(_07645_),
    .B1(_07906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08046_));
 sky130_fd_sc_hd__a21oi_2 _17179_ (.A1(_07812_),
    .A2(_07906_),
    .B1(_08045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08047_));
 sky130_fd_sc_hd__a21o_2 _17180_ (.A1(_07812_),
    .A2(_07906_),
    .B1(_08045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08048_));
 sky130_fd_sc_hd__a2bb2o_2 _17181_ (.A1_N(_07642_),
    .A2_N(_07811_),
    .B1(_08043_),
    .B2(_08044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08049_));
 sky130_fd_sc_hd__and3_2 _17182_ (.A(_07812_),
    .B(_07906_),
    .C(_08045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08050_));
 sky130_fd_sc_hd__nand2_2 _17183_ (.A(\a_l[11] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_2 _17184_ (.A(\a_l[13] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08052_));
 sky130_fd_sc_hd__a22oi_2 _17185_ (.A1(\a_l[13] ),
    .A2(\b_h[6] ),
    .B1(\b_h[7] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08053_));
 sky130_fd_sc_hd__nand2_2 _17186_ (.A(_07925_),
    .B(_08052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08054_));
 sky130_fd_sc_hd__nand2_2 _17187_ (.A(\a_l[13] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08055_));
 sky130_fd_sc_hd__and4_2 _17188_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08056_));
 sky130_fd_sc_hd__nand4_2 _17189_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08057_));
 sky130_fd_sc_hd__o2111ai_2 _17190_ (.A1(_07923_),
    .A2(_08055_),
    .B1(\a_l[11] ),
    .C1(\b_h[8] ),
    .D1(_08054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08058_));
 sky130_fd_sc_hd__o2bb2ai_2 _17191_ (.A1_N(_08054_),
    .A2_N(_08057_),
    .B1(_09297_),
    .B2(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08059_));
 sky130_fd_sc_hd__a21oi_2 _17192_ (.A1(_08054_),
    .A2(_08057_),
    .B1(_08051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08060_));
 sky130_fd_sc_hd__a21o_2 _17193_ (.A1(_08054_),
    .A2(_08057_),
    .B1(_08051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08061_));
 sky130_fd_sc_hd__nand2_2 _17194_ (.A(_08051_),
    .B(_08057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08062_));
 sky130_fd_sc_hd__nand3_2 _17195_ (.A(_08059_),
    .B(_07902_),
    .C(_08058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08063_));
 sky130_fd_sc_hd__a31oi_2 _17196_ (.A1(_08051_),
    .A2(_08054_),
    .A3(_08057_),
    .B1(_07902_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08064_));
 sky130_fd_sc_hd__o21ai_2 _17197_ (.A1(_08053_),
    .A2(_08062_),
    .B1(_07903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_2 _17198_ (.A(_08064_),
    .B(_08061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08066_));
 sky130_fd_sc_hd__o21a_2 _17199_ (.A1(_08060_),
    .A2(_08065_),
    .B1(_08063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08067_));
 sky130_fd_sc_hd__o21ai_2 _17200_ (.A1(_08060_),
    .A2(_08065_),
    .B1(_08063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08068_));
 sky130_fd_sc_hd__o21ai_2 _17201_ (.A1(_07921_),
    .A2(_07926_),
    .B1(_07924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08069_));
 sky130_fd_sc_hd__a31o_2 _17202_ (.A1(\a_l[10] ),
    .A2(_07924_),
    .A3(\b_h[8] ),
    .B1(_07926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08070_));
 sky130_fd_sc_hd__o211ai_2 _17203_ (.A1(_08060_),
    .A2(_08065_),
    .B1(_08069_),
    .C1(_08063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08071_));
 sky130_fd_sc_hd__nand2_2 _17204_ (.A(_08068_),
    .B(_08070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08072_));
 sky130_fd_sc_hd__o211ai_2 _17205_ (.A1(_08047_),
    .A2(_08050_),
    .B1(_08071_),
    .C1(_08072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08073_));
 sky130_fd_sc_hd__a21oi_2 _17206_ (.A1(_08063_),
    .A2(_08066_),
    .B1(_08070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08074_));
 sky130_fd_sc_hd__o211ai_2 _17207_ (.A1(_08060_),
    .A2(_08065_),
    .B1(_08070_),
    .C1(_08063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08075_));
 sky130_fd_sc_hd__o211a_2 _17208_ (.A1(_08049_),
    .A2(_07907_),
    .B1(_08048_),
    .C1(_08075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08076_));
 sky130_fd_sc_hd__o211ai_2 _17209_ (.A1(_08049_),
    .A2(_07907_),
    .B1(_08048_),
    .C1(_08075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08077_));
 sky130_fd_sc_hd__o21ai_2 _17210_ (.A1(_08067_),
    .A2(_08070_),
    .B1(_08076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08078_));
 sky130_fd_sc_hd__o21ai_2 _17211_ (.A1(_08074_),
    .A2(_08077_),
    .B1(_08073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08079_));
 sky130_fd_sc_hd__o211ai_2 _17212_ (.A1(_07912_),
    .A2(_07898_),
    .B1(_07939_),
    .C1(_07937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08080_));
 sky130_fd_sc_hd__o21ai_2 _17213_ (.A1(_07936_),
    .A2(_07941_),
    .B1(_07916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08081_));
 sky130_fd_sc_hd__o21a_2 _17214_ (.A1(_07936_),
    .A2(_07941_),
    .B1(_07916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08082_));
 sky130_fd_sc_hd__a21oi_2 _17215_ (.A1(_07916_),
    .A2(_08080_),
    .B1(_08079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08083_));
 sky130_fd_sc_hd__nand3_2 _17216_ (.A(_08081_),
    .B(_08078_),
    .C(_08073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08084_));
 sky130_fd_sc_hd__a21oi_2 _17217_ (.A1(_08073_),
    .A2(_08078_),
    .B1(_08081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08085_));
 sky130_fd_sc_hd__nand2_2 _17218_ (.A(_08079_),
    .B(_08082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08086_));
 sky130_fd_sc_hd__o31a_2 _17219_ (.A1(_07958_),
    .A2(_07960_),
    .A3(_07950_),
    .B1(_07974_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08087_));
 sky130_fd_sc_hd__o21ai_2 _17220_ (.A1(_07971_),
    .A2(_07972_),
    .B1(_07964_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08088_));
 sky130_fd_sc_hd__o211a_2 _17221_ (.A1(_07967_),
    .A2(_07970_),
    .B1(_07973_),
    .C1(_07963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08089_));
 sky130_fd_sc_hd__a21o_2 _17222_ (.A1(_07963_),
    .A2(_07975_),
    .B1(_07965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08090_));
 sky130_fd_sc_hd__nand2_2 _17223_ (.A(_07963_),
    .B(_08088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08091_));
 sky130_fd_sc_hd__o2bb2ai_2 _17224_ (.A1_N(_07920_),
    .A2_N(_07935_),
    .B1(_07933_),
    .B2(_07928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08092_));
 sky130_fd_sc_hd__a21boi_2 _17225_ (.A1(_07920_),
    .A2(_07935_),
    .B1_N(_07934_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08093_));
 sky130_fd_sc_hd__nand2_2 _17226_ (.A(\a_l[5] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08094_));
 sky130_fd_sc_hd__a22oi_2 _17227_ (.A1(\a_l[7] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08095_));
 sky130_fd_sc_hd__and4_2 _17228_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08096_));
 sky130_fd_sc_hd__nand4_2 _17229_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08097_));
 sky130_fd_sc_hd__o21bai_2 _17230_ (.A1(_08095_),
    .A2(_08096_),
    .B1_N(_08094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08098_));
 sky130_fd_sc_hd__o21a_2 _17231_ (.A1(_09210_),
    .A2(_09668_),
    .B1(_08097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08099_));
 sky130_fd_sc_hd__o21ai_2 _17232_ (.A1(_09210_),
    .A2(_09668_),
    .B1(_08097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08100_));
 sky130_fd_sc_hd__o21ai_2 _17233_ (.A1(_08095_),
    .A2(_08100_),
    .B1(_08098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08101_));
 sky130_fd_sc_hd__o2bb2ai_2 _17234_ (.A1_N(_07951_),
    .A2_N(_07954_),
    .B1(_02338_),
    .B2(_06985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08102_));
 sky130_fd_sc_hd__a21boi_2 _17235_ (.A1(_07954_),
    .A2(_07951_),
    .B1_N(_07955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08103_));
 sky130_fd_sc_hd__nand2_2 _17236_ (.A(\a_l[8] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08104_));
 sky130_fd_sc_hd__nand2_2 _17237_ (.A(\a_l[9] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08105_));
 sky130_fd_sc_hd__nand2_2 _17238_ (.A(\a_l[10] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08106_));
 sky130_fd_sc_hd__a22oi_2 _17239_ (.A1(\a_l[10] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08107_));
 sky130_fd_sc_hd__nand2_2 _17240_ (.A(_08105_),
    .B(_08106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08108_));
 sky130_fd_sc_hd__nand4_2 _17241_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08109_));
 sky130_fd_sc_hd__nand2_2 _17242_ (.A(_08104_),
    .B(_08109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08110_));
 sky130_fd_sc_hd__a21o_2 _17243_ (.A1(_08108_),
    .A2(_08109_),
    .B1(_08104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08111_));
 sky130_fd_sc_hd__o2bb2ai_2 _17244_ (.A1_N(_08108_),
    .A2_N(_08109_),
    .B1(_09253_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08112_));
 sky130_fd_sc_hd__o2111ai_2 _17245_ (.A1(_02338_),
    .A2(_07100_),
    .B1(\a_l[8] ),
    .C1(\b_h[11] ),
    .D1(_08108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08113_));
 sky130_fd_sc_hd__o211ai_2 _17246_ (.A1(_08110_),
    .A2(_08107_),
    .B1(_08103_),
    .C1(_08111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08114_));
 sky130_fd_sc_hd__inv_2 _17247_ (.A(_08114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08115_));
 sky130_fd_sc_hd__nand3_2 _17248_ (.A(_08112_),
    .B(_08113_),
    .C(_08102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08116_));
 sky130_fd_sc_hd__nand2_2 _17249_ (.A(_08114_),
    .B(_08116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08117_));
 sky130_fd_sc_hd__nand2_2 _17250_ (.A(_08117_),
    .B(_08101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08118_));
 sky130_fd_sc_hd__o211a_2 _17251_ (.A1(_08100_),
    .A2(_08095_),
    .B1(_08098_),
    .C1(_08116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08119_));
 sky130_fd_sc_hd__o2111ai_2 _17252_ (.A1(_08100_),
    .A2(_08095_),
    .B1(_08098_),
    .C1(_08114_),
    .D1(_08116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08120_));
 sky130_fd_sc_hd__nand3_2 _17253_ (.A(_08114_),
    .B(_08116_),
    .C(_08101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08121_));
 sky130_fd_sc_hd__a21o_2 _17254_ (.A1(_08114_),
    .A2(_08116_),
    .B1(_08101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08122_));
 sky130_fd_sc_hd__nand3_2 _17255_ (.A(_08122_),
    .B(_08092_),
    .C(_08121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08123_));
 sky130_fd_sc_hd__nand3_2 _17256_ (.A(_08093_),
    .B(_08118_),
    .C(_08120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08124_));
 sky130_fd_sc_hd__a31oi_2 _17257_ (.A1(_08122_),
    .A2(_08092_),
    .A3(_08121_),
    .B1(_08091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08125_));
 sky130_fd_sc_hd__nand2_2 _17258_ (.A(_08124_),
    .B(_08090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08126_));
 sky130_fd_sc_hd__o211a_2 _17259_ (.A1(_07965_),
    .A2(_08089_),
    .B1(_08123_),
    .C1(_08124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08127_));
 sky130_fd_sc_hd__nand2_2 _17260_ (.A(_08125_),
    .B(_08124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08128_));
 sky130_fd_sc_hd__a2bb2oi_2 _17261_ (.A1_N(_07962_),
    .A2_N(_08087_),
    .B1(_08123_),
    .B2(_08124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08129_));
 sky130_fd_sc_hd__a22o_2 _17262_ (.A1(_07963_),
    .A2(_08088_),
    .B1(_08123_),
    .B2(_08124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08130_));
 sky130_fd_sc_hd__a21oi_2 _17263_ (.A1(_08124_),
    .A2(_08125_),
    .B1(_08129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08131_));
 sky130_fd_sc_hd__o211ai_2 _17264_ (.A1(_08127_),
    .A2(_08129_),
    .B1(_08084_),
    .C1(_08086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08132_));
 sky130_fd_sc_hd__o21ai_2 _17265_ (.A1(_08083_),
    .A2(_08085_),
    .B1(_08131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08133_));
 sky130_fd_sc_hd__o2bb2ai_2 _17266_ (.A1_N(_08084_),
    .A2_N(_08086_),
    .B1(_08127_),
    .B2(_08129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08134_));
 sky130_fd_sc_hd__a22oi_2 _17267_ (.A1(_08125_),
    .A2(_08124_),
    .B1(_08082_),
    .B2(_08079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08135_));
 sky130_fd_sc_hd__nand3_2 _17268_ (.A(_08086_),
    .B(_08128_),
    .C(_08130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08136_));
 sky130_fd_sc_hd__nand4_2 _17269_ (.A(_08084_),
    .B(_08086_),
    .C(_08128_),
    .D(_08130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08137_));
 sky130_fd_sc_hd__o211ai_2 _17270_ (.A1(_08083_),
    .A2(_08136_),
    .B1(_08134_),
    .C1(_07992_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08138_));
 sky130_fd_sc_hd__nand3_2 _17271_ (.A(_07993_),
    .B(_08132_),
    .C(_08133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08139_));
 sky130_fd_sc_hd__and3_2 _17272_ (.A(_08138_),
    .B(_08139_),
    .C(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08140_));
 sky130_fd_sc_hd__nand3_2 _17273_ (.A(_08138_),
    .B(_08139_),
    .C(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08141_));
 sky130_fd_sc_hd__a21oi_2 _17274_ (.A1(_08138_),
    .A2(_08139_),
    .B1(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08142_));
 sky130_fd_sc_hd__a21o_2 _17275_ (.A1(_08138_),
    .A2(_08139_),
    .B1(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08143_));
 sky130_fd_sc_hd__a2bb2oi_2 _17276_ (.A1_N(_08000_),
    .A2_N(_08031_),
    .B1(_08141_),
    .B2(_08143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08144_));
 sky130_fd_sc_hd__o22ai_2 _17277_ (.A1(_08000_),
    .A2(_08031_),
    .B1(_08140_),
    .B2(_08142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08145_));
 sky130_fd_sc_hd__o21ai_2 _17278_ (.A1(_07998_),
    .A2(_08003_),
    .B1(_08143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08146_));
 sky130_fd_sc_hd__o211ai_2 _17279_ (.A1(_07998_),
    .A2(_08003_),
    .B1(_08141_),
    .C1(_08143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08147_));
 sky130_fd_sc_hd__nand2_2 _17280_ (.A(_08145_),
    .B(_08147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08148_));
 sky130_fd_sc_hd__a21oi_2 _17281_ (.A1(_07892_),
    .A2(_07887_),
    .B1(_07890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08149_));
 sky130_fd_sc_hd__inv_2 _17282_ (.A(_08149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08150_));
 sky130_fd_sc_hd__and3_2 _17283_ (.A(_08145_),
    .B(_08147_),
    .C(_08150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08151_));
 sky130_fd_sc_hd__nand2_2 _17284_ (.A(_08148_),
    .B(_08150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08152_));
 sky130_fd_sc_hd__o211ai_2 _17285_ (.A1(_08140_),
    .A2(_08146_),
    .B1(_08149_),
    .C1(_08145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08153_));
 sky130_fd_sc_hd__a31oi_2 _17286_ (.A1(_08004_),
    .A2(_08005_),
    .A3(_08007_),
    .B1(_08013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08154_));
 sky130_fd_sc_hd__a31oi_2 _17287_ (.A1(_08006_),
    .A2(_08002_),
    .A3(_08001_),
    .B1(_08014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08155_));
 sky130_fd_sc_hd__o211ai_2 _17288_ (.A1(_08008_),
    .A2(_08154_),
    .B1(_08153_),
    .C1(_08152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08156_));
 sky130_fd_sc_hd__o2bb2ai_2 _17289_ (.A1_N(_08149_),
    .A2_N(_08148_),
    .B1(_08010_),
    .B2(_08155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08157_));
 sky130_fd_sc_hd__o2bb2ai_2 _17290_ (.A1_N(_08152_),
    .A2_N(_08153_),
    .B1(_08155_),
    .B2(_08010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08158_));
 sky130_fd_sc_hd__o21a_2 _17291_ (.A1(_08151_),
    .A2(_08157_),
    .B1(_08156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08159_));
 sky130_fd_sc_hd__o21ai_2 _17292_ (.A1(_08151_),
    .A2(_08157_),
    .B1(_08156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08160_));
 sky130_fd_sc_hd__a21oi_2 _17293_ (.A1(_08020_),
    .A2(_08030_),
    .B1(_08160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08161_));
 sky130_fd_sc_hd__a31o_2 _17294_ (.A1(_08020_),
    .A2(_08030_),
    .A3(_08160_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08162_));
 sky130_fd_sc_hd__nor2_2 _17295_ (.A(_08161_),
    .B(_08162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00357_));
 sky130_fd_sc_hd__o22ai_2 _17296_ (.A1(_08140_),
    .A2(_08146_),
    .B1(_08149_),
    .B2(_08144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08163_));
 sky130_fd_sc_hd__a32oi_2 _17297_ (.A1(_07992_),
    .A2(_08134_),
    .A3(_08137_),
    .B1(_08139_),
    .B2(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08164_));
 sky130_fd_sc_hd__a32o_2 _17298_ (.A1(_07992_),
    .A2(_08134_),
    .A3(_08137_),
    .B1(_08139_),
    .B2(_08040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08165_));
 sky130_fd_sc_hd__o21ai_2 _17299_ (.A1(_08104_),
    .A2(_08107_),
    .B1(_08109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08166_));
 sky130_fd_sc_hd__nand2_2 _17300_ (.A(_08108_),
    .B(_08110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_2 _17301_ (.A(\a_l[9] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08168_));
 sky130_fd_sc_hd__a22oi_2 _17302_ (.A1(\a_l[11] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08169_));
 sky130_fd_sc_hd__nor2_2 _17303_ (.A(_02338_),
    .B(_07234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08170_));
 sky130_fd_sc_hd__nand4_2 _17304_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08171_));
 sky130_fd_sc_hd__o21ai_2 _17305_ (.A1(_08169_),
    .A2(_08170_),
    .B1(_08168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08172_));
 sky130_fd_sc_hd__a41o_2 _17306_ (.A1(\a_l[10] ),
    .A2(\a_l[11] ),
    .A3(\b_h[9] ),
    .A4(\b_h[10] ),
    .B1(_08168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08173_));
 sky130_fd_sc_hd__o21ai_2 _17307_ (.A1(_02338_),
    .A2(_07234_),
    .B1(_08168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08174_));
 sky130_fd_sc_hd__o21bai_2 _17308_ (.A1(_08169_),
    .A2(_08170_),
    .B1_N(_08168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08175_));
 sky130_fd_sc_hd__o211a_2 _17309_ (.A1(_08174_),
    .A2(_08169_),
    .B1(_08167_),
    .C1(_08175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08176_));
 sky130_fd_sc_hd__o211ai_2 _17310_ (.A1(_08174_),
    .A2(_08169_),
    .B1(_08167_),
    .C1(_08175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08177_));
 sky130_fd_sc_hd__o211ai_2 _17311_ (.A1(_08169_),
    .A2(_08173_),
    .B1(_08166_),
    .C1(_08172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08178_));
 sky130_fd_sc_hd__inv_2 _17312_ (.A(_08178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08179_));
 sky130_fd_sc_hd__and4_2 _17313_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08180_));
 sky130_fd_sc_hd__a22oi_2 _17314_ (.A1(\a_l[8] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08181_));
 sky130_fd_sc_hd__a22o_2 _17315_ (.A1(\a_l[8] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08182_));
 sky130_fd_sc_hd__o2111a_2 _17316_ (.A1(_02589_),
    .A2(_06867_),
    .B1(\a_l[6] ),
    .C1(\b_h[14] ),
    .D1(_08182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08183_));
 sky130_fd_sc_hd__o2111ai_2 _17317_ (.A1(_02589_),
    .A2(_06867_),
    .B1(\a_l[6] ),
    .C1(\b_h[14] ),
    .D1(_08182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08184_));
 sky130_fd_sc_hd__o22a_2 _17318_ (.A1(_09231_),
    .A2(_09668_),
    .B1(_08180_),
    .B2(_08181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08185_));
 sky130_fd_sc_hd__o22ai_2 _17319_ (.A1(_09231_),
    .A2(_09668_),
    .B1(_08180_),
    .B2(_08181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08186_));
 sky130_fd_sc_hd__o2bb2ai_2 _17320_ (.A1_N(_08177_),
    .A2_N(_08178_),
    .B1(_08183_),
    .B2(_08185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08187_));
 sky130_fd_sc_hd__nand3_2 _17321_ (.A(_08178_),
    .B(_08184_),
    .C(_08186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08188_));
 sky130_fd_sc_hd__nand4_2 _17322_ (.A(_08177_),
    .B(_08178_),
    .C(_08184_),
    .D(_08186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08189_));
 sky130_fd_sc_hd__inv_2 _17323_ (.A(_08189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08190_));
 sky130_fd_sc_hd__a22oi_2 _17324_ (.A1(_08061_),
    .A2(_08064_),
    .B1(_08063_),
    .B2(_08069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08191_));
 sky130_fd_sc_hd__a21oi_2 _17325_ (.A1(_08187_),
    .A2(_08189_),
    .B1(_08191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08192_));
 sky130_fd_sc_hd__a21o_2 _17326_ (.A1(_08187_),
    .A2(_08189_),
    .B1(_08191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08193_));
 sky130_fd_sc_hd__o211a_2 _17327_ (.A1(_08176_),
    .A2(_08188_),
    .B1(_08191_),
    .C1(_08187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08194_));
 sky130_fd_sc_hd__nand3_2 _17328_ (.A(_08187_),
    .B(_08189_),
    .C(_08191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08195_));
 sky130_fd_sc_hd__nand2_2 _17329_ (.A(_08114_),
    .B(_08101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08196_));
 sky130_fd_sc_hd__nand2_2 _17330_ (.A(_08116_),
    .B(_08196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08197_));
 sky130_fd_sc_hd__o22a_2 _17331_ (.A1(_08115_),
    .A2(_08119_),
    .B1(_08192_),
    .B2(_08194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08198_));
 sky130_fd_sc_hd__o22ai_2 _17332_ (.A1(_08115_),
    .A2(_08119_),
    .B1(_08192_),
    .B2(_08194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08199_));
 sky130_fd_sc_hd__nand3_2 _17333_ (.A(_08193_),
    .B(_08195_),
    .C(_08197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08200_));
 sky130_fd_sc_hd__o21ai_2 _17334_ (.A1(_08192_),
    .A2(_08194_),
    .B1(_08197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08201_));
 sky130_fd_sc_hd__o211ai_2 _17335_ (.A1(_08115_),
    .A2(_08119_),
    .B1(_08193_),
    .C1(_08195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08202_));
 sky130_fd_sc_hd__o22ai_2 _17336_ (.A1(_08045_),
    .A2(_08046_),
    .B1(_08074_),
    .B2(_08077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08203_));
 sky130_fd_sc_hd__and3_2 _17337_ (.A(_08054_),
    .B(\b_h[8] ),
    .C(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08204_));
 sky130_fd_sc_hd__a31o_2 _17338_ (.A1(\a_l[11] ),
    .A2(_08054_),
    .A3(\b_h[8] ),
    .B1(_08056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08205_));
 sky130_fd_sc_hd__and2_2 _17339_ (.A(\a_l[12] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08206_));
 sky130_fd_sc_hd__nand2_2 _17340_ (.A(\a_l[14] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08207_));
 sky130_fd_sc_hd__nand2_2 _17341_ (.A(_08055_),
    .B(_08207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08208_));
 sky130_fd_sc_hd__and2_2 _17342_ (.A(\a_l[14] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08209_));
 sky130_fd_sc_hd__nand2_2 _17343_ (.A(\a_l[14] ),
    .B(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08210_));
 sky130_fd_sc_hd__o2bb2ai_2 _17344_ (.A1_N(_08055_),
    .A2_N(_08207_),
    .B1(_08210_),
    .B2(_08052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08211_));
 sky130_fd_sc_hd__o221ai_2 _17345_ (.A1(_09319_),
    .A2(_09613_),
    .B1(_08052_),
    .B2(_08210_),
    .C1(_08208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_2 _17346_ (.A(_08211_),
    .B(_08206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08213_));
 sky130_fd_sc_hd__o211a_2 _17347_ (.A1(_08052_),
    .A2(_08210_),
    .B1(_08206_),
    .C1(_08208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08214_));
 sky130_fd_sc_hd__o211ai_2 _17348_ (.A1(_08052_),
    .A2(_08210_),
    .B1(_08206_),
    .C1(_08208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08215_));
 sky130_fd_sc_hd__o21ai_2 _17349_ (.A1(_09319_),
    .A2(_09613_),
    .B1(_08211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08216_));
 sky130_fd_sc_hd__nand2_2 _17350_ (.A(_08215_),
    .B(_08216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_2 _17351_ (.A(_08216_),
    .B(_08042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08218_));
 sky130_fd_sc_hd__nand3_2 _17352_ (.A(_08216_),
    .B(_08042_),
    .C(_08215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08219_));
 sky130_fd_sc_hd__nand3_2 _17353_ (.A(_08043_),
    .B(_08212_),
    .C(_08213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08220_));
 sky130_fd_sc_hd__a21oi_2 _17354_ (.A1(_08219_),
    .A2(_08220_),
    .B1(_08205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08221_));
 sky130_fd_sc_hd__a22o_2 _17355_ (.A1(_08054_),
    .A2(_08062_),
    .B1(_08219_),
    .B2(_08220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08222_));
 sky130_fd_sc_hd__o211ai_2 _17356_ (.A1(_08056_),
    .A2(_08204_),
    .B1(_08219_),
    .C1(_08220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08223_));
 sky130_fd_sc_hd__nand3b_2 _17357_ (.A_N(_08205_),
    .B(_08219_),
    .C(_08220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08224_));
 sky130_fd_sc_hd__a21oi_2 _17358_ (.A1(_08217_),
    .A2(_08205_),
    .B1(_08041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08225_));
 sky130_fd_sc_hd__nand2_2 _17359_ (.A(_08225_),
    .B(_08224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08226_));
 sky130_fd_sc_hd__nand2_2 _17360_ (.A(_08223_),
    .B(_08041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08227_));
 sky130_fd_sc_hd__nand4_2 _17361_ (.A(_08222_),
    .B(_08223_),
    .C(\a_l[15] ),
    .D(\b_h[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08228_));
 sky130_fd_sc_hd__o21ai_2 _17362_ (.A1(_08221_),
    .A2(_08227_),
    .B1(_08226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08229_));
 sky130_fd_sc_hd__o211ai_2 _17363_ (.A1(_08077_),
    .A2(_08074_),
    .B1(_08048_),
    .C1(_08229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08230_));
 sky130_fd_sc_hd__inv_2 _17364_ (.A(_08230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08231_));
 sky130_fd_sc_hd__nand3_2 _17365_ (.A(_08203_),
    .B(_08226_),
    .C(_08228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_2 _17366_ (.A(_08230_),
    .B(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08233_));
 sky130_fd_sc_hd__a21boi_2 _17367_ (.A1(_08199_),
    .A2(_08200_),
    .B1_N(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08234_));
 sky130_fd_sc_hd__nand3_2 _17368_ (.A(_08201_),
    .B(_08202_),
    .C(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08235_));
 sky130_fd_sc_hd__nand4_2 _17369_ (.A(_08201_),
    .B(_08202_),
    .C(_08230_),
    .D(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08236_));
 sky130_fd_sc_hd__nand3_2 _17370_ (.A(_08199_),
    .B(_08200_),
    .C(_08233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08237_));
 sky130_fd_sc_hd__a21oi_2 _17371_ (.A1(_08135_),
    .A2(_08130_),
    .B1(_08083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08238_));
 sky130_fd_sc_hd__o21ai_2 _17372_ (.A1(_08079_),
    .A2(_08082_),
    .B1(_08136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08239_));
 sky130_fd_sc_hd__nand3_2 _17373_ (.A(_08238_),
    .B(_08237_),
    .C(_08236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08240_));
 sky130_fd_sc_hd__a22o_2 _17374_ (.A1(_08199_),
    .A2(_08200_),
    .B1(_08230_),
    .B2(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08241_));
 sky130_fd_sc_hd__nand3_2 _17375_ (.A(_08200_),
    .B(_08230_),
    .C(_08232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08242_));
 sky130_fd_sc_hd__a2bb2oi_2 _17376_ (.A1_N(_08198_),
    .A2_N(_08242_),
    .B1(_08084_),
    .B2(_08136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08243_));
 sky130_fd_sc_hd__o211ai_2 _17377_ (.A1(_08198_),
    .A2(_08242_),
    .B1(_08241_),
    .C1(_08239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08244_));
 sky130_fd_sc_hd__a21oi_2 _17378_ (.A1(_08094_),
    .A2(_08097_),
    .B1(_08095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08245_));
 sky130_fd_sc_hd__o21ai_2 _17379_ (.A1(_07962_),
    .A2(_08087_),
    .B1(_08123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08246_));
 sky130_fd_sc_hd__nand3_2 _17380_ (.A(_08124_),
    .B(_08245_),
    .C(_08246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08247_));
 sky130_fd_sc_hd__o211ai_2 _17381_ (.A1(_08095_),
    .A2(_08099_),
    .B1(_08123_),
    .C1(_08126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08248_));
 sky130_fd_sc_hd__inv_2 _17382_ (.A(_08248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08249_));
 sky130_fd_sc_hd__nand2_2 _17383_ (.A(_08247_),
    .B(_08248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08250_));
 sky130_fd_sc_hd__nor2_2 _17384_ (.A(_09210_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_2 _17385_ (.A(\a_l[5] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08252_));
 sky130_fd_sc_hd__a31o_2 _17386_ (.A1(_08124_),
    .A2(_08245_),
    .A3(_08246_),
    .B1(_08251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08253_));
 sky130_fd_sc_hd__and3_2 _17387_ (.A(_08247_),
    .B(_08248_),
    .C(_08252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08254_));
 sky130_fd_sc_hd__and3_2 _17388_ (.A(_08250_),
    .B(\b_h[15] ),
    .C(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08255_));
 sky130_fd_sc_hd__nand2_2 _17389_ (.A(_08250_),
    .B(_08251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08256_));
 sky130_fd_sc_hd__o2bb2a_2 _17390_ (.A1_N(_08247_),
    .A2_N(_08248_),
    .B1(_09210_),
    .B2(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08257_));
 sky130_fd_sc_hd__and3_2 _17391_ (.A(_08247_),
    .B(_08248_),
    .C(_08251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08258_));
 sky130_fd_sc_hd__o21ai_2 _17392_ (.A1(_08249_),
    .A2(_08253_),
    .B1(_08256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08259_));
 sky130_fd_sc_hd__nand3b_2 _17393_ (.A_N(_08259_),
    .B(_08244_),
    .C(_08240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08260_));
 sky130_fd_sc_hd__o2bb2ai_2 _17394_ (.A1_N(_08240_),
    .A2_N(_08244_),
    .B1(_08254_),
    .B2(_08255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08261_));
 sky130_fd_sc_hd__o211ai_2 _17395_ (.A1(_08254_),
    .A2(_08255_),
    .B1(_08240_),
    .C1(_08244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08262_));
 sky130_fd_sc_hd__o2bb2ai_2 _17396_ (.A1_N(_08240_),
    .A2_N(_08244_),
    .B1(_08257_),
    .B2(_08258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08263_));
 sky130_fd_sc_hd__nand3_2 _17397_ (.A(_08165_),
    .B(_08262_),
    .C(_08263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08264_));
 sky130_fd_sc_hd__nand3_2 _17398_ (.A(_08261_),
    .B(_08164_),
    .C(_08260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08265_));
 sky130_fd_sc_hd__nand2_2 _17399_ (.A(_08036_),
    .B(_08038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08266_));
 sky130_fd_sc_hd__a21bo_2 _17400_ (.A1(_08264_),
    .A2(_08265_),
    .B1_N(_08266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08267_));
 sky130_fd_sc_hd__nand4_2 _17401_ (.A(_08036_),
    .B(_08038_),
    .C(_08264_),
    .D(_08265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08268_));
 sky130_fd_sc_hd__a21o_2 _17402_ (.A1(_08267_),
    .A2(_08268_),
    .B1(_08163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08269_));
 sky130_fd_sc_hd__nand3_2 _17403_ (.A(_08163_),
    .B(_08267_),
    .C(_08268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08270_));
 sky130_fd_sc_hd__nand2_2 _17404_ (.A(_08269_),
    .B(_08270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08271_));
 sky130_fd_sc_hd__o21ai_2 _17405_ (.A1(_08017_),
    .A2(_08019_),
    .B1(_08158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08272_));
 sky130_fd_sc_hd__nand2_2 _17406_ (.A(_08156_),
    .B(_08272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08273_));
 sky130_fd_sc_hd__nor2_2 _17407_ (.A(_08023_),
    .B(_08160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08274_));
 sky130_fd_sc_hd__nand4_2 _17408_ (.A(_08020_),
    .B(_08021_),
    .C(_08156_),
    .D(_08158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08275_));
 sky130_fd_sc_hd__nor2_2 _17409_ (.A(_08025_),
    .B(_08275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08276_));
 sky130_fd_sc_hd__nand4_2 _17410_ (.A(_07584_),
    .B(_08024_),
    .C(_08274_),
    .D(_07586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08277_));
 sky130_fd_sc_hd__nand4_2 _17411_ (.A(_08022_),
    .B(_08159_),
    .C(_08026_),
    .D(_07879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08278_));
 sky130_fd_sc_hd__a22oi_2 _17412_ (.A1(_08156_),
    .A2(_08272_),
    .B1(_08274_),
    .B2(_08027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08279_));
 sky130_fd_sc_hd__nand2_2 _17413_ (.A(_08277_),
    .B(_08279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08280_));
 sky130_fd_sc_hd__a21o_2 _17414_ (.A1(_08269_),
    .A2(_08270_),
    .B1(_08280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08281_));
 sky130_fd_sc_hd__a31o_2 _17415_ (.A1(_08277_),
    .A2(_08278_),
    .A3(_08273_),
    .B1(_08271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08282_));
 sky130_fd_sc_hd__and3_2 _17416_ (.A(_09690_),
    .B(_08281_),
    .C(_08282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00358_));
 sky130_fd_sc_hd__a22o_2 _17417_ (.A1(_08243_),
    .A2(_08241_),
    .B1(_08240_),
    .B2(_08259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08283_));
 sky130_fd_sc_hd__a22oi_2 _17418_ (.A1(_08243_),
    .A2(_08241_),
    .B1(_08240_),
    .B2(_08259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08284_));
 sky130_fd_sc_hd__nand2_2 _17419_ (.A(_08230_),
    .B(_08235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08285_));
 sky130_fd_sc_hd__nand2_2 _17420_ (.A(\a_l[15] ),
    .B(\b_h[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08286_));
 sky130_fd_sc_hd__nand4_2 _17421_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[6] ),
    .D(\b_h[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_2 _17422_ (.A(_08210_),
    .B(_08286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08288_));
 sky130_fd_sc_hd__a22o_2 _17423_ (.A1(\a_l[13] ),
    .A2(\b_h[8] ),
    .B1(_08287_),
    .B2(_08288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08289_));
 sky130_fd_sc_hd__nand4_2 _17424_ (.A(_08288_),
    .B(\b_h[8] ),
    .C(\a_l[13] ),
    .D(_08287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08290_));
 sky130_fd_sc_hd__a2bb2o_2 _17425_ (.A1_N(_08052_),
    .A2_N(_08210_),
    .B1(_08206_),
    .B2(_08208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08291_));
 sky130_fd_sc_hd__a21o_2 _17426_ (.A1(_08289_),
    .A2(_08290_),
    .B1(_08291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08292_));
 sky130_fd_sc_hd__and3_2 _17427_ (.A(_08289_),
    .B(_08291_),
    .C(_08290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08293_));
 sky130_fd_sc_hd__nand3_2 _17428_ (.A(_08289_),
    .B(_08291_),
    .C(_08290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08294_));
 sky130_fd_sc_hd__nand2_2 _17429_ (.A(_08292_),
    .B(_08294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08295_));
 sky130_fd_sc_hd__nand3_2 _17430_ (.A(_08222_),
    .B(_08292_),
    .C(_08294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08296_));
 sky130_fd_sc_hd__nor3_2 _17431_ (.A(_08295_),
    .B(_08221_),
    .C(_08227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08297_));
 sky130_fd_sc_hd__o2bb2a_2 _17432_ (.A1_N(_08292_),
    .A2_N(_08294_),
    .B1(_08221_),
    .B2(_08227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08298_));
 sky130_fd_sc_hd__o21ai_2 _17433_ (.A1(_08221_),
    .A2(_08227_),
    .B1(_08295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08299_));
 sky130_fd_sc_hd__o21a_2 _17434_ (.A1(_08227_),
    .A2(_08296_),
    .B1(_08299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08300_));
 sky130_fd_sc_hd__o21a_2 _17435_ (.A1(_08176_),
    .A2(_08188_),
    .B1(_08178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08301_));
 sky130_fd_sc_hd__a21o_2 _17436_ (.A1(_08168_),
    .A2(_08171_),
    .B1(_08169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08302_));
 sky130_fd_sc_hd__a21oi_2 _17437_ (.A1(_08168_),
    .A2(_08171_),
    .B1(_08169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08303_));
 sky130_fd_sc_hd__nand2_2 _17438_ (.A(\a_l[10] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_2 _17439_ (.A(\a_l[11] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_2 _17440_ (.A(\a_l[12] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08306_));
 sky130_fd_sc_hd__a22oi_2 _17441_ (.A1(\a_l[12] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_2 _17442_ (.A(_08305_),
    .B(_08306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08308_));
 sky130_fd_sc_hd__nand2_2 _17443_ (.A(\a_l[12] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08309_));
 sky130_fd_sc_hd__nand4_2 _17444_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08310_));
 sky130_fd_sc_hd__nand3_2 _17445_ (.A(_08310_),
    .B(\b_h[11] ),
    .C(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08311_));
 sky130_fd_sc_hd__o2bb2ai_2 _17446_ (.A1_N(_08308_),
    .A2_N(_08310_),
    .B1(_09286_),
    .B2(_09646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08312_));
 sky130_fd_sc_hd__o211ai_2 _17447_ (.A1(_08311_),
    .A2(_08307_),
    .B1(_08303_),
    .C1(_08312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08313_));
 sky130_fd_sc_hd__o21ai_2 _17448_ (.A1(_08305_),
    .A2(_08306_),
    .B1(_08304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08314_));
 sky130_fd_sc_hd__a21o_2 _17449_ (.A1(_08308_),
    .A2(_08310_),
    .B1(_08304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08315_));
 sky130_fd_sc_hd__o211a_2 _17450_ (.A1(_08307_),
    .A2(_08314_),
    .B1(_08302_),
    .C1(_08315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08316_));
 sky130_fd_sc_hd__o211ai_2 _17451_ (.A1(_08307_),
    .A2(_08314_),
    .B1(_08302_),
    .C1(_08315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08317_));
 sky130_fd_sc_hd__a22o_2 _17452_ (.A1(\a_l[9] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08318_));
 sky130_fd_sc_hd__o21ai_2 _17453_ (.A1(_02589_),
    .A2(_06985_),
    .B1(_08318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08319_));
 sky130_fd_sc_hd__o2111a_2 _17454_ (.A1(_02589_),
    .A2(_06985_),
    .B1(\a_l[7] ),
    .C1(\b_h[14] ),
    .D1(_08318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08320_));
 sky130_fd_sc_hd__o2111ai_2 _17455_ (.A1(_02589_),
    .A2(_06985_),
    .B1(\a_l[7] ),
    .C1(\b_h[14] ),
    .D1(_08318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08321_));
 sky130_fd_sc_hd__o21a_2 _17456_ (.A1(_09242_),
    .A2(_09668_),
    .B1(_08319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08322_));
 sky130_fd_sc_hd__o21ai_2 _17457_ (.A1(_09242_),
    .A2(_09668_),
    .B1(_08319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08323_));
 sky130_fd_sc_hd__o2bb2ai_2 _17458_ (.A1_N(_08313_),
    .A2_N(_08317_),
    .B1(_08320_),
    .B2(_08322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08324_));
 sky130_fd_sc_hd__nand3_2 _17459_ (.A(_08313_),
    .B(_08321_),
    .C(_08323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08325_));
 sky130_fd_sc_hd__nand4_2 _17460_ (.A(_08313_),
    .B(_08317_),
    .C(_08321_),
    .D(_08323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08326_));
 sky130_fd_sc_hd__o2bb2ai_2 _17461_ (.A1_N(_08205_),
    .A2_N(_08220_),
    .B1(_08218_),
    .B2(_08214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08327_));
 sky130_fd_sc_hd__a21oi_2 _17462_ (.A1(_08324_),
    .A2(_08326_),
    .B1(_08327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08328_));
 sky130_fd_sc_hd__a21o_2 _17463_ (.A1(_08324_),
    .A2(_08326_),
    .B1(_08327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08329_));
 sky130_fd_sc_hd__o211a_2 _17464_ (.A1(_08316_),
    .A2(_08325_),
    .B1(_08327_),
    .C1(_08324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08330_));
 sky130_fd_sc_hd__o211ai_2 _17465_ (.A1(_08316_),
    .A2(_08325_),
    .B1(_08327_),
    .C1(_08324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08331_));
 sky130_fd_sc_hd__o211ai_2 _17466_ (.A1(_08179_),
    .A2(_08190_),
    .B1(_08329_),
    .C1(_08331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08332_));
 sky130_fd_sc_hd__o21ai_2 _17467_ (.A1(_08328_),
    .A2(_08330_),
    .B1(_08301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08333_));
 sky130_fd_sc_hd__nand3_2 _17468_ (.A(_08329_),
    .B(_08331_),
    .C(_08301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08334_));
 sky130_fd_sc_hd__o22ai_2 _17469_ (.A1(_08179_),
    .A2(_08190_),
    .B1(_08328_),
    .B2(_08330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08335_));
 sky130_fd_sc_hd__and3_2 _17470_ (.A(_08333_),
    .B(_08300_),
    .C(_08332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08336_));
 sky130_fd_sc_hd__nand3_2 _17471_ (.A(_08333_),
    .B(_08300_),
    .C(_08332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08337_));
 sky130_fd_sc_hd__o211ai_2 _17472_ (.A1(_08297_),
    .A2(_08298_),
    .B1(_08334_),
    .C1(_08335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08338_));
 sky130_fd_sc_hd__nand2_2 _17473_ (.A(_08337_),
    .B(_08338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08339_));
 sky130_fd_sc_hd__nand3_2 _17474_ (.A(_08230_),
    .B(_08235_),
    .C(_08338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08340_));
 sky130_fd_sc_hd__and4_2 _17475_ (.A(_08230_),
    .B(_08235_),
    .C(_08337_),
    .D(_08338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08341_));
 sky130_fd_sc_hd__nor2_2 _17476_ (.A(_09231_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08342_));
 sky130_fd_sc_hd__a31o_2 _17477_ (.A1(_08182_),
    .A2(\b_h[14] ),
    .A3(\a_l[6] ),
    .B1(_08180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08343_));
 sky130_fd_sc_hd__a31oi_2 _17478_ (.A1(_08187_),
    .A2(_08189_),
    .A3(_08191_),
    .B1(_08197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08344_));
 sky130_fd_sc_hd__o21ai_2 _17479_ (.A1(_08115_),
    .A2(_08119_),
    .B1(_08195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08345_));
 sky130_fd_sc_hd__o21bai_2 _17480_ (.A1(_08192_),
    .A2(_08344_),
    .B1_N(_08343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08346_));
 sky130_fd_sc_hd__o211ai_2 _17481_ (.A1(_08180_),
    .A2(_08183_),
    .B1(_08193_),
    .C1(_08345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08347_));
 sky130_fd_sc_hd__and3_2 _17482_ (.A(_08346_),
    .B(_08347_),
    .C(_08342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08348_));
 sky130_fd_sc_hd__a21oi_2 _17483_ (.A1(_08346_),
    .A2(_08347_),
    .B1(_08342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08349_));
 sky130_fd_sc_hd__nor2_2 _17484_ (.A(_08348_),
    .B(_08349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08350_));
 sky130_fd_sc_hd__o21ai_2 _17485_ (.A1(_08231_),
    .A2(_08234_),
    .B1(_08339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08351_));
 sky130_fd_sc_hd__a21oi_2 _17486_ (.A1(_08350_),
    .A2(_08351_),
    .B1(_08341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08352_));
 sky130_fd_sc_hd__a2bb2o_2 _17487_ (.A1_N(_08336_),
    .A2_N(_08340_),
    .B1(_08351_),
    .B2(_08350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08353_));
 sky130_fd_sc_hd__o21ai_2 _17488_ (.A1(_08336_),
    .A2(_08340_),
    .B1(_08351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08354_));
 sky130_fd_sc_hd__o211ai_2 _17489_ (.A1(_08336_),
    .A2(_08340_),
    .B1(_08351_),
    .C1(_08350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08355_));
 sky130_fd_sc_hd__o21ai_2 _17490_ (.A1(_08348_),
    .A2(_08349_),
    .B1(_08354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08356_));
 sky130_fd_sc_hd__o2bb2ai_2 _17491_ (.A1_N(_08285_),
    .A2_N(_08339_),
    .B1(_08348_),
    .B2(_08349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08357_));
 sky130_fd_sc_hd__nand2_2 _17492_ (.A(_08354_),
    .B(_08350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08358_));
 sky130_fd_sc_hd__nand3_2 _17493_ (.A(_08283_),
    .B(_08355_),
    .C(_08356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08359_));
 sky130_fd_sc_hd__o211ai_2 _17494_ (.A1(_08357_),
    .A2(_08341_),
    .B1(_08284_),
    .C1(_08358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08360_));
 sky130_fd_sc_hd__o21ai_2 _17495_ (.A1(_08252_),
    .A2(_08249_),
    .B1(_08247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08361_));
 sky130_fd_sc_hd__a22o_2 _17496_ (.A1(_08248_),
    .A2(_08253_),
    .B1(_08359_),
    .B2(_08360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08362_));
 sky130_fd_sc_hd__nand4_2 _17497_ (.A(_08248_),
    .B(_08253_),
    .C(_08359_),
    .D(_08360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08363_));
 sky130_fd_sc_hd__a21boi_2 _17498_ (.A1(_08264_),
    .A2(_08266_),
    .B1_N(_08265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08364_));
 sky130_fd_sc_hd__a21oi_2 _17499_ (.A1(_08362_),
    .A2(_08363_),
    .B1(_08364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08365_));
 sky130_fd_sc_hd__a21o_2 _17500_ (.A1(_08362_),
    .A2(_08363_),
    .B1(_08364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08366_));
 sky130_fd_sc_hd__nand3_2 _17501_ (.A(_08362_),
    .B(_08363_),
    .C(_08364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08367_));
 sky130_fd_sc_hd__nand2_2 _17502_ (.A(_08366_),
    .B(_08367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08368_));
 sky130_fd_sc_hd__a21oi_2 _17503_ (.A1(_08270_),
    .A2(_08282_),
    .B1(_08368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08369_));
 sky130_fd_sc_hd__and3_2 _17504_ (.A(_08270_),
    .B(_08282_),
    .C(_08368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08370_));
 sky130_fd_sc_hd__nor3_2 _17505_ (.A(rst),
    .B(_08369_),
    .C(_08370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_2 _17506_ (.A(_08360_),
    .B(_08361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08371_));
 sky130_fd_sc_hd__nand2_2 _17507_ (.A(_08359_),
    .B(_08371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08372_));
 sky130_fd_sc_hd__a21bo_2 _17508_ (.A1(_08342_),
    .A2(_08346_),
    .B1_N(_08347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08373_));
 sky130_fd_sc_hd__o211ai_2 _17509_ (.A1(_08228_),
    .A2(_08295_),
    .B1(_08334_),
    .C1(_08335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08374_));
 sky130_fd_sc_hd__nor2_2 _17510_ (.A(_09373_),
    .B(_09613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08375_));
 sky130_fd_sc_hd__nand2_2 _17511_ (.A(\a_l[15] ),
    .B(\b_h[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08376_));
 sky130_fd_sc_hd__and3_2 _17512_ (.A(\a_l[15] ),
    .B(\b_h[8] ),
    .C(_08209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08377_));
 sky130_fd_sc_hd__a22oi_2 _17513_ (.A1(\a_l[15] ),
    .A2(\b_h[7] ),
    .B1(\b_h[8] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08378_));
 sky130_fd_sc_hd__o221a_2 _17514_ (.A1(_08210_),
    .A2(_08286_),
    .B1(_08377_),
    .B2(_08378_),
    .C1(_08290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08379_));
 sky130_fd_sc_hd__a221oi_2 _17515_ (.A1(_08209_),
    .A2(_08375_),
    .B1(_08290_),
    .B2(_08287_),
    .C1(_08378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08380_));
 sky130_fd_sc_hd__a221o_2 _17516_ (.A1(_08209_),
    .A2(_08375_),
    .B1(_08290_),
    .B2(_08287_),
    .C1(_08378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08381_));
 sky130_fd_sc_hd__or2_2 _17517_ (.A(_08379_),
    .B(_08380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08382_));
 sky130_fd_sc_hd__inv_2 _17518_ (.A(_08382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08383_));
 sky130_fd_sc_hd__and2_2 _17519_ (.A(\a_l[8] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08384_));
 sky130_fd_sc_hd__nand2_2 _17520_ (.A(\a_l[9] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08385_));
 sky130_fd_sc_hd__a22o_2 _17521_ (.A1(\a_l[10] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08386_));
 sky130_fd_sc_hd__a21o_2 _17522_ (.A1(\a_l[10] ),
    .A2(\b_h[12] ),
    .B1(_08385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08387_));
 sky130_fd_sc_hd__o211a_2 _17523_ (.A1(_02589_),
    .A2(_07100_),
    .B1(_08384_),
    .C1(_08386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08388_));
 sky130_fd_sc_hd__a31oi_2 _17524_ (.A1(\a_l[10] ),
    .A2(\b_h[12] ),
    .A3(_08385_),
    .B1(_08384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08389_));
 sky130_fd_sc_hd__a21oi_2 _17525_ (.A1(_08387_),
    .A2(_08389_),
    .B1(_08388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08390_));
 sky130_fd_sc_hd__a21o_2 _17526_ (.A1(_08387_),
    .A2(_08389_),
    .B1(_08388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08391_));
 sky130_fd_sc_hd__a21o_2 _17527_ (.A1(_08304_),
    .A2(_08310_),
    .B1(_08307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08392_));
 sky130_fd_sc_hd__a21oi_2 _17528_ (.A1(_08304_),
    .A2(_08310_),
    .B1(_08307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08393_));
 sky130_fd_sc_hd__nand2_2 _17529_ (.A(\a_l[11] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08394_));
 sky130_fd_sc_hd__nand2_2 _17530_ (.A(\a_l[13] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08395_));
 sky130_fd_sc_hd__a22oi_2 _17531_ (.A1(\a_l[13] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08396_));
 sky130_fd_sc_hd__nand2_2 _17532_ (.A(_08309_),
    .B(_08395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08397_));
 sky130_fd_sc_hd__and4_2 _17533_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08398_));
 sky130_fd_sc_hd__nand4_2 _17534_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08399_));
 sky130_fd_sc_hd__nand3_2 _17535_ (.A(_08399_),
    .B(\b_h[11] ),
    .C(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08400_));
 sky130_fd_sc_hd__o22ai_2 _17536_ (.A1(_09297_),
    .A2(_09646_),
    .B1(_08396_),
    .B2(_08398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08401_));
 sky130_fd_sc_hd__o22a_2 _17537_ (.A1(_09297_),
    .A2(_09646_),
    .B1(_08309_),
    .B2(_08395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08402_));
 sky130_fd_sc_hd__o211ai_2 _17538_ (.A1(_09297_),
    .A2(_09646_),
    .B1(_08397_),
    .C1(_08399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08403_));
 sky130_fd_sc_hd__a21o_2 _17539_ (.A1(_08397_),
    .A2(_08399_),
    .B1(_08394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08404_));
 sky130_fd_sc_hd__o211ai_2 _17540_ (.A1(_08400_),
    .A2(_08396_),
    .B1(_08393_),
    .C1(_08401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08405_));
 sky130_fd_sc_hd__and3_2 _17541_ (.A(_08404_),
    .B(_08392_),
    .C(_08403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08406_));
 sky130_fd_sc_hd__nand3_2 _17542_ (.A(_08404_),
    .B(_08392_),
    .C(_08403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_2 _17543_ (.A(_08405_),
    .B(_08407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08408_));
 sky130_fd_sc_hd__nand3_2 _17544_ (.A(_08391_),
    .B(_08405_),
    .C(_08407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08409_));
 sky130_fd_sc_hd__nand2_2 _17545_ (.A(_08408_),
    .B(_08390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08410_));
 sky130_fd_sc_hd__a21o_2 _17546_ (.A1(_08405_),
    .A2(_08407_),
    .B1(_08390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08411_));
 sky130_fd_sc_hd__nand3_2 _17547_ (.A(_08390_),
    .B(_08405_),
    .C(_08407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08412_));
 sky130_fd_sc_hd__nand3_2 _17548_ (.A(_08294_),
    .B(_08409_),
    .C(_08410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08413_));
 sky130_fd_sc_hd__and3_2 _17549_ (.A(_08411_),
    .B(_08412_),
    .C(_08293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08414_));
 sky130_fd_sc_hd__nand3_2 _17550_ (.A(_08411_),
    .B(_08412_),
    .C(_08293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08415_));
 sky130_fd_sc_hd__nand2_2 _17551_ (.A(_08413_),
    .B(_08415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08416_));
 sky130_fd_sc_hd__o21a_2 _17552_ (.A1(_08316_),
    .A2(_08325_),
    .B1(_08313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08417_));
 sky130_fd_sc_hd__o21ai_2 _17553_ (.A1(_08316_),
    .A2(_08325_),
    .B1(_08313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_2 _17554_ (.A(_08416_),
    .B(_08418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_2 _17555_ (.A(_08413_),
    .B(_08417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08420_));
 sky130_fd_sc_hd__nand4_2 _17556_ (.A(_08313_),
    .B(_08326_),
    .C(_08413_),
    .D(_08415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08421_));
 sky130_fd_sc_hd__nand3_2 _17557_ (.A(_08413_),
    .B(_08415_),
    .C(_08418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08422_));
 sky130_fd_sc_hd__a21o_2 _17558_ (.A1(_08413_),
    .A2(_08415_),
    .B1(_08418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08423_));
 sky130_fd_sc_hd__o21a_2 _17559_ (.A1(_08414_),
    .A2(_08420_),
    .B1(_08419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08424_));
 sky130_fd_sc_hd__a21oi_2 _17560_ (.A1(_08419_),
    .A2(_08421_),
    .B1(_08382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08425_));
 sky130_fd_sc_hd__nand3_2 _17561_ (.A(_08423_),
    .B(_08383_),
    .C(_08422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08426_));
 sky130_fd_sc_hd__o211a_2 _17562_ (.A1(_08420_),
    .A2(_08414_),
    .B1(_08382_),
    .C1(_08419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08427_));
 sky130_fd_sc_hd__o211ai_2 _17563_ (.A1(_08420_),
    .A2(_08414_),
    .B1(_08382_),
    .C1(_08419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08428_));
 sky130_fd_sc_hd__nand4_2 _17564_ (.A(_08299_),
    .B(_08374_),
    .C(_08426_),
    .D(_08428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08429_));
 sky130_fd_sc_hd__a22oi_2 _17565_ (.A1(_08299_),
    .A2(_08374_),
    .B1(_08426_),
    .B2(_08428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08430_));
 sky130_fd_sc_hd__o2bb2ai_2 _17566_ (.A1_N(_08299_),
    .A2_N(_08374_),
    .B1(_08425_),
    .B2(_08427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08431_));
 sky130_fd_sc_hd__nor2_2 _17567_ (.A(_09242_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08432_));
 sky130_fd_sc_hd__o31a_2 _17568_ (.A1(_09253_),
    .A2(_09275_),
    .A3(_02589_),
    .B1(_08321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08433_));
 sky130_fd_sc_hd__a31o_2 _17569_ (.A1(\a_l[8] ),
    .A2(\a_l[9] ),
    .A3(_02588_),
    .B1(_08320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08434_));
 sky130_fd_sc_hd__nand2_2 _17570_ (.A(_08331_),
    .B(_08301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08435_));
 sky130_fd_sc_hd__nand3_2 _17571_ (.A(_08329_),
    .B(_08434_),
    .C(_08435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08436_));
 sky130_fd_sc_hd__o211ai_2 _17572_ (.A1(_08301_),
    .A2(_08328_),
    .B1(_08331_),
    .C1(_08433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08437_));
 sky130_fd_sc_hd__a21oi_2 _17573_ (.A1(_08436_),
    .A2(_08437_),
    .B1(_08432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08438_));
 sky130_fd_sc_hd__a22o_2 _17574_ (.A1(\a_l[7] ),
    .A2(\b_h[15] ),
    .B1(_08436_),
    .B2(_08437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08439_));
 sky130_fd_sc_hd__and3_2 _17575_ (.A(_08436_),
    .B(_08437_),
    .C(_08432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08440_));
 sky130_fd_sc_hd__nand4_2 _17576_ (.A(_08437_),
    .B(\a_l[7] ),
    .C(_08436_),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08441_));
 sky130_fd_sc_hd__nor2_2 _17577_ (.A(_08438_),
    .B(_08440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08442_));
 sky130_fd_sc_hd__nand2_2 _17578_ (.A(_08439_),
    .B(_08441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08443_));
 sky130_fd_sc_hd__o211ai_2 _17579_ (.A1(_08438_),
    .A2(_08440_),
    .B1(_08429_),
    .C1(_08431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08444_));
 sky130_fd_sc_hd__a21o_2 _17580_ (.A1(_08429_),
    .A2(_08431_),
    .B1(_08443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08445_));
 sky130_fd_sc_hd__a21o_2 _17581_ (.A1(_08429_),
    .A2(_08431_),
    .B1(_08442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08446_));
 sky130_fd_sc_hd__nand4_2 _17582_ (.A(_08429_),
    .B(_08431_),
    .C(_08439_),
    .D(_08441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08447_));
 sky130_fd_sc_hd__nand3_2 _17583_ (.A(_08353_),
    .B(_08446_),
    .C(_08447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08448_));
 sky130_fd_sc_hd__and3_2 _17584_ (.A(_08445_),
    .B(_08352_),
    .C(_08444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08449_));
 sky130_fd_sc_hd__nand3_2 _17585_ (.A(_08445_),
    .B(_08352_),
    .C(_08444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08450_));
 sky130_fd_sc_hd__a21oi_2 _17586_ (.A1(_08448_),
    .A2(_08450_),
    .B1(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08451_));
 sky130_fd_sc_hd__a21o_2 _17587_ (.A1(_08448_),
    .A2(_08450_),
    .B1(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08452_));
 sky130_fd_sc_hd__nand2_2 _17588_ (.A(_08450_),
    .B(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08453_));
 sky130_fd_sc_hd__and3_2 _17589_ (.A(_08448_),
    .B(_08450_),
    .C(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08454_));
 sky130_fd_sc_hd__nand3_2 _17590_ (.A(_08448_),
    .B(_08450_),
    .C(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08455_));
 sky130_fd_sc_hd__o21bai_2 _17591_ (.A1(_08451_),
    .A2(_08454_),
    .B1_N(_08372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08456_));
 sky130_fd_sc_hd__nand3_2 _17592_ (.A(_08452_),
    .B(_08455_),
    .C(_08372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08457_));
 sky130_fd_sc_hd__nand2_2 _17593_ (.A(_08456_),
    .B(_08457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08458_));
 sky130_fd_sc_hd__a21o_2 _17594_ (.A1(_08270_),
    .A2(_08367_),
    .B1(_08365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08459_));
 sky130_fd_sc_hd__a21oi_2 _17595_ (.A1(_08270_),
    .A2(_08367_),
    .B1(_08365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08460_));
 sky130_fd_sc_hd__and4_2 _17596_ (.A(_08269_),
    .B(_08270_),
    .C(_08366_),
    .D(_08367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08461_));
 sky130_fd_sc_hd__a21oi_2 _17597_ (.A1(_08280_),
    .A2(_08461_),
    .B1(_08460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08462_));
 sky130_fd_sc_hd__nor2_2 _17598_ (.A(_08458_),
    .B(_08462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08463_));
 sky130_fd_sc_hd__o21ai_2 _17599_ (.A1(_08458_),
    .A2(_08462_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08464_));
 sky130_fd_sc_hd__a21oi_2 _17600_ (.A1(_08458_),
    .A2(_08462_),
    .B1(_08464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00360_));
 sky130_fd_sc_hd__a31oi_2 _17601_ (.A1(_08353_),
    .A2(_08446_),
    .A3(_08447_),
    .B1(_08373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08465_));
 sky130_fd_sc_hd__nand2_2 _17602_ (.A(_08448_),
    .B(_08453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08466_));
 sky130_fd_sc_hd__a31o_2 _17603_ (.A1(\a_l[9] ),
    .A2(\a_l[10] ),
    .A3(_02588_),
    .B1(_08388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08467_));
 sky130_fd_sc_hd__nand2_2 _17604_ (.A(_08415_),
    .B(_08417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08468_));
 sky130_fd_sc_hd__nand2_2 _17605_ (.A(_08413_),
    .B(_08418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08469_));
 sky130_fd_sc_hd__nand3_2 _17606_ (.A(_08413_),
    .B(_08467_),
    .C(_08468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08470_));
 sky130_fd_sc_hd__nand3b_2 _17607_ (.A_N(_08467_),
    .B(_08469_),
    .C(_08415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08471_));
 sky130_fd_sc_hd__nor2_2 _17608_ (.A(_09253_),
    .B(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08472_));
 sky130_fd_sc_hd__a31o_2 _17609_ (.A1(_08413_),
    .A2(_08467_),
    .A3(_08468_),
    .B1(_08472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08473_));
 sky130_fd_sc_hd__a21oi_2 _17610_ (.A1(_08470_),
    .A2(_08471_),
    .B1(_08472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08474_));
 sky130_fd_sc_hd__a21o_2 _17611_ (.A1(_08470_),
    .A2(_08471_),
    .B1(_08472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08475_));
 sky130_fd_sc_hd__and3_2 _17612_ (.A(_08470_),
    .B(_08471_),
    .C(_08472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08476_));
 sky130_fd_sc_hd__nand4_2 _17613_ (.A(_08470_),
    .B(_08471_),
    .C(\a_l[8] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08477_));
 sky130_fd_sc_hd__nand2_2 _17614_ (.A(_08475_),
    .B(_08477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08478_));
 sky130_fd_sc_hd__and3_2 _17615_ (.A(_08210_),
    .B(\b_h[8] ),
    .C(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08479_));
 sky130_fd_sc_hd__nand2_2 _17616_ (.A(\a_l[10] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_2 _17617_ (.A(\a_l[11] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08481_));
 sky130_fd_sc_hd__and3_2 _17618_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(_02588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08482_));
 sky130_fd_sc_hd__nand4_2 _17619_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08483_));
 sky130_fd_sc_hd__nand2_2 _17620_ (.A(_08480_),
    .B(_08481_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08484_));
 sky130_fd_sc_hd__and4_2 _17621_ (.A(_08484_),
    .B(\b_h[14] ),
    .C(\a_l[9] ),
    .D(_08483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08485_));
 sky130_fd_sc_hd__o2111ai_2 _17622_ (.A1(_02589_),
    .A2(_07234_),
    .B1(\a_l[9] ),
    .C1(\b_h[14] ),
    .D1(_08484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08486_));
 sky130_fd_sc_hd__a22o_2 _17623_ (.A1(\a_l[9] ),
    .A2(\b_h[14] ),
    .B1(_08483_),
    .B2(_08484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08487_));
 sky130_fd_sc_hd__nand2_2 _17624_ (.A(_08486_),
    .B(_08487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08488_));
 sky130_fd_sc_hd__a21oi_2 _17625_ (.A1(_08309_),
    .A2(_08395_),
    .B1(_08394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08489_));
 sky130_fd_sc_hd__nand2_2 _17626_ (.A(\a_l[13] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_2 _17627_ (.A(\a_l[14] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08491_));
 sky130_fd_sc_hd__a22oi_2 _17628_ (.A1(\a_l[14] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08492_));
 sky130_fd_sc_hd__nand2_2 _17629_ (.A(_08490_),
    .B(_08491_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08493_));
 sky130_fd_sc_hd__nand2_2 _17630_ (.A(\a_l[14] ),
    .B(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08494_));
 sky130_fd_sc_hd__nand4_2 _17631_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08495_));
 sky130_fd_sc_hd__o2bb2ai_2 _17632_ (.A1_N(_08490_),
    .A2_N(_08491_),
    .B1(_08494_),
    .B2(_08395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08496_));
 sky130_fd_sc_hd__nand2_2 _17633_ (.A(\a_l[12] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08497_));
 sky130_fd_sc_hd__o2111ai_2 _17634_ (.A1(_08395_),
    .A2(_08494_),
    .B1(\a_l[12] ),
    .C1(\b_h[11] ),
    .D1(_08493_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08498_));
 sky130_fd_sc_hd__nand2_2 _17635_ (.A(_08496_),
    .B(_08497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08499_));
 sky130_fd_sc_hd__nand2_2 _17636_ (.A(_08498_),
    .B(_08499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08500_));
 sky130_fd_sc_hd__o211a_2 _17637_ (.A1(_08398_),
    .A2(_08489_),
    .B1(_08498_),
    .C1(_08499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08501_));
 sky130_fd_sc_hd__o211ai_2 _17638_ (.A1(_08398_),
    .A2(_08489_),
    .B1(_08498_),
    .C1(_08499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08502_));
 sky130_fd_sc_hd__a2bb2oi_2 _17639_ (.A1_N(_08396_),
    .A2_N(_08402_),
    .B1(_08498_),
    .B2(_08499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08503_));
 sky130_fd_sc_hd__o21ai_2 _17640_ (.A1(_08396_),
    .A2(_08402_),
    .B1(_08500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08504_));
 sky130_fd_sc_hd__nand3_2 _17641_ (.A(_08488_),
    .B(_08502_),
    .C(_08504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08505_));
 sky130_fd_sc_hd__o21bai_2 _17642_ (.A1(_08501_),
    .A2(_08503_),
    .B1_N(_08488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08506_));
 sky130_fd_sc_hd__and4_2 _17643_ (.A(_08486_),
    .B(_08487_),
    .C(_08502_),
    .D(_08504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08507_));
 sky130_fd_sc_hd__nand3b_2 _17644_ (.A_N(_08488_),
    .B(_08502_),
    .C(_08504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08508_));
 sky130_fd_sc_hd__o21ai_2 _17645_ (.A1(_08501_),
    .A2(_08503_),
    .B1(_08488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08509_));
 sky130_fd_sc_hd__nand2_2 _17646_ (.A(_08509_),
    .B(_08380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08510_));
 sky130_fd_sc_hd__nand3_2 _17647_ (.A(_08509_),
    .B(_08380_),
    .C(_08508_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08511_));
 sky130_fd_sc_hd__nand3_2 _17648_ (.A(_08381_),
    .B(_08505_),
    .C(_08506_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08512_));
 sky130_fd_sc_hd__nand2_2 _17649_ (.A(_08511_),
    .B(_08512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08513_));
 sky130_fd_sc_hd__and2_2 _17650_ (.A(_08391_),
    .B(_08405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08514_));
 sky130_fd_sc_hd__o21ai_2 _17651_ (.A1(_08391_),
    .A2(_08406_),
    .B1(_08405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08515_));
 sky130_fd_sc_hd__a31o_2 _17652_ (.A1(_08392_),
    .A2(_08403_),
    .A3(_08404_),
    .B1(_08514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08516_));
 sky130_fd_sc_hd__nand3_2 _17653_ (.A(_08511_),
    .B(_08512_),
    .C(_08515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08517_));
 sky130_fd_sc_hd__o2bb2ai_2 _17654_ (.A1_N(_08511_),
    .A2_N(_08512_),
    .B1(_08514_),
    .B2(_08406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08518_));
 sky130_fd_sc_hd__a21boi_2 _17655_ (.A1(_08513_),
    .A2(_08516_),
    .B1_N(_08479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08519_));
 sky130_fd_sc_hd__nand4_2 _17656_ (.A(_08210_),
    .B(_08518_),
    .C(_08375_),
    .D(_08517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08520_));
 sky130_fd_sc_hd__a22oi_2 _17657_ (.A1(_08375_),
    .A2(_08210_),
    .B1(_08518_),
    .B2(_08517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08521_));
 sky130_fd_sc_hd__o2bb2ai_2 _17658_ (.A1_N(_08517_),
    .A2_N(_08518_),
    .B1(_08209_),
    .B2(_08376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08522_));
 sky130_fd_sc_hd__a211oi_2 _17659_ (.A1(_08519_),
    .A2(_08517_),
    .B1(_08426_),
    .C1(_08521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08523_));
 sky130_fd_sc_hd__nand3_2 _17660_ (.A(_08522_),
    .B(_08425_),
    .C(_08520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08524_));
 sky130_fd_sc_hd__a21oi_2 _17661_ (.A1(_08520_),
    .A2(_08522_),
    .B1(_08425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08525_));
 sky130_fd_sc_hd__o2bb2ai_2 _17662_ (.A1_N(_08520_),
    .A2_N(_08522_),
    .B1(_08382_),
    .B2(_08424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08526_));
 sky130_fd_sc_hd__a21o_2 _17663_ (.A1(_08524_),
    .A2(_08526_),
    .B1(_08478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08527_));
 sky130_fd_sc_hd__o211ai_2 _17664_ (.A1(_08474_),
    .A2(_08476_),
    .B1(_08524_),
    .C1(_08526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08528_));
 sky130_fd_sc_hd__o21ai_2 _17665_ (.A1(_08523_),
    .A2(_08525_),
    .B1(_08478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08529_));
 sky130_fd_sc_hd__nand4_2 _17666_ (.A(_08475_),
    .B(_08477_),
    .C(_08524_),
    .D(_08526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08530_));
 sky130_fd_sc_hd__o21ai_2 _17667_ (.A1(_08443_),
    .A2(_08430_),
    .B1(_08429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08531_));
 sky130_fd_sc_hd__a21boi_2 _17668_ (.A1(_08442_),
    .A2(_08431_),
    .B1_N(_08429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08532_));
 sky130_fd_sc_hd__nand3_2 _17669_ (.A(_08527_),
    .B(_08528_),
    .C(_08532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08533_));
 sky130_fd_sc_hd__nand3_2 _17670_ (.A(_08529_),
    .B(_08530_),
    .C(_08531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08534_));
 sky130_fd_sc_hd__a21bo_2 _17671_ (.A1(_08432_),
    .A2(_08437_),
    .B1_N(_08436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08535_));
 sky130_fd_sc_hd__inv_2 _17672_ (.A(_08535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08536_));
 sky130_fd_sc_hd__nand3_2 _17673_ (.A(_08533_),
    .B(_08534_),
    .C(_08535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08537_));
 sky130_fd_sc_hd__a21o_2 _17674_ (.A1(_08533_),
    .A2(_08534_),
    .B1(_08535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08538_));
 sky130_fd_sc_hd__nand3_2 _17675_ (.A(_08533_),
    .B(_08534_),
    .C(_08536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08539_));
 sky130_fd_sc_hd__a21o_2 _17676_ (.A1(_08533_),
    .A2(_08534_),
    .B1(_08536_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08540_));
 sky130_fd_sc_hd__o211ai_2 _17677_ (.A1(_08449_),
    .A2(_08465_),
    .B1(_08539_),
    .C1(_08540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08541_));
 sky130_fd_sc_hd__nand3_2 _17678_ (.A(_08538_),
    .B(_08466_),
    .C(_08537_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08542_));
 sky130_fd_sc_hd__and2_2 _17679_ (.A(_08541_),
    .B(_08542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08543_));
 sky130_fd_sc_hd__o21ai_2 _17680_ (.A1(_08458_),
    .A2(_08462_),
    .B1(_08457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08544_));
 sky130_fd_sc_hd__a31o_2 _17681_ (.A1(_08372_),
    .A2(_08452_),
    .A3(_08455_),
    .B1(_08543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08545_));
 sky130_fd_sc_hd__nand2_2 _17682_ (.A(_08544_),
    .B(_08543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08546_));
 sky130_fd_sc_hd__o211a_2 _17683_ (.A1(_08545_),
    .A2(_08463_),
    .B1(_09690_),
    .C1(_08546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00361_));
 sky130_fd_sc_hd__o21ai_2 _17684_ (.A1(_08474_),
    .A2(_08476_),
    .B1(_08524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08547_));
 sky130_fd_sc_hd__o21ai_2 _17685_ (.A1(_08478_),
    .A2(_08525_),
    .B1(_08524_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08548_));
 sky130_fd_sc_hd__nand2_2 _17686_ (.A(_08526_),
    .B(_08547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08549_));
 sky130_fd_sc_hd__nand2_2 _17687_ (.A(\a_l[11] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_2 _17688_ (.A(\a_l[12] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_2 _17689_ (.A(_08550_),
    .B(_08551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_2 _17690_ (.A(\a_l[12] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08553_));
 sky130_fd_sc_hd__and4_2 _17691_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08554_));
 sky130_fd_sc_hd__nand4_2 _17692_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08555_));
 sky130_fd_sc_hd__and2_2 _17693_ (.A(\a_l[10] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08556_));
 sky130_fd_sc_hd__and3_2 _17694_ (.A(_08552_),
    .B(_08556_),
    .C(_08555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08557_));
 sky130_fd_sc_hd__o2111ai_2 _17695_ (.A1(_08481_),
    .A2(_08553_),
    .B1(\a_l[10] ),
    .C1(\b_h[14] ),
    .D1(_08552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08558_));
 sky130_fd_sc_hd__a21oi_2 _17696_ (.A1(_08552_),
    .A2(_08555_),
    .B1(_08556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08559_));
 sky130_fd_sc_hd__a22o_2 _17697_ (.A1(\a_l[10] ),
    .A2(\b_h[14] ),
    .B1(_08552_),
    .B2(_08555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08560_));
 sky130_fd_sc_hd__nor2_2 _17698_ (.A(_08557_),
    .B(_08559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08561_));
 sky130_fd_sc_hd__nand2_2 _17699_ (.A(_08558_),
    .B(_08560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08562_));
 sky130_fd_sc_hd__nand2_2 _17700_ (.A(\a_l[13] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08563_));
 sky130_fd_sc_hd__nand4_2 _17701_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[9] ),
    .D(\b_h[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08564_));
 sky130_fd_sc_hd__nand2_2 _17702_ (.A(\a_l[15] ),
    .B(\b_h[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08565_));
 sky130_fd_sc_hd__a22oi_2 _17703_ (.A1(\a_l[15] ),
    .A2(\b_h[9] ),
    .B1(\b_h[10] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08566_));
 sky130_fd_sc_hd__nand2_2 _17704_ (.A(_08494_),
    .B(_08565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08567_));
 sky130_fd_sc_hd__a2bb2oi_2 _17705_ (.A1_N(_09340_),
    .A2_N(_09646_),
    .B1(_08564_),
    .B2(_08567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08568_));
 sky130_fd_sc_hd__a22o_2 _17706_ (.A1(\a_l[13] ),
    .A2(\b_h[11] ),
    .B1(_08564_),
    .B2(_08567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08569_));
 sky130_fd_sc_hd__nand3_2 _17707_ (.A(_08564_),
    .B(\b_h[11] ),
    .C(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08570_));
 sky130_fd_sc_hd__nor2_2 _17708_ (.A(_08566_),
    .B(_08570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08571_));
 sky130_fd_sc_hd__nand4_2 _17709_ (.A(_08567_),
    .B(\b_h[11] ),
    .C(\a_l[13] ),
    .D(_08564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08572_));
 sky130_fd_sc_hd__o21ai_2 _17710_ (.A1(_08497_),
    .A2(_08492_),
    .B1(_08495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08573_));
 sky130_fd_sc_hd__a21oi_2 _17711_ (.A1(_08569_),
    .A2(_08572_),
    .B1(_08573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08574_));
 sky130_fd_sc_hd__o21bai_2 _17712_ (.A1(_08568_),
    .A2(_08571_),
    .B1_N(_08573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08575_));
 sky130_fd_sc_hd__nand3_2 _17713_ (.A(_08569_),
    .B(_08572_),
    .C(_08573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08576_));
 sky130_fd_sc_hd__a21oi_2 _17714_ (.A1(_08575_),
    .A2(_08576_),
    .B1(_08561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08577_));
 sky130_fd_sc_hd__a21o_2 _17715_ (.A1(_08575_),
    .A2(_08576_),
    .B1(_08561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08578_));
 sky130_fd_sc_hd__nand3_2 _17716_ (.A(_08561_),
    .B(_08575_),
    .C(_08576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08579_));
 sky130_fd_sc_hd__a21oi_2 _17717_ (.A1(_08575_),
    .A2(_08576_),
    .B1(_08562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08580_));
 sky130_fd_sc_hd__a21o_2 _17718_ (.A1(_08575_),
    .A2(_08576_),
    .B1(_08562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08581_));
 sky130_fd_sc_hd__a31oi_2 _17719_ (.A1(_08562_),
    .A2(_08575_),
    .A3(_08576_),
    .B1(_08377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08582_));
 sky130_fd_sc_hd__a31o_2 _17720_ (.A1(_08562_),
    .A2(_08575_),
    .A3(_08576_),
    .B1(_08377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08583_));
 sky130_fd_sc_hd__nand2_2 _17721_ (.A(_08582_),
    .B(_08581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_2 _17722_ (.A(_08579_),
    .B(_08377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08585_));
 sky130_fd_sc_hd__nand4_2 _17723_ (.A(_08578_),
    .B(_08579_),
    .C(_08209_),
    .D(_08375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08586_));
 sky130_fd_sc_hd__o21ai_2 _17724_ (.A1(_08488_),
    .A2(_08503_),
    .B1(_08502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08587_));
 sky130_fd_sc_hd__o221ai_2 _17725_ (.A1(_08577_),
    .A2(_08585_),
    .B1(_08580_),
    .B2(_08583_),
    .C1(_08587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08588_));
 sky130_fd_sc_hd__a21o_2 _17726_ (.A1(_08584_),
    .A2(_08586_),
    .B1(_08587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08589_));
 sky130_fd_sc_hd__nand2_2 _17727_ (.A(_08588_),
    .B(_08589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08590_));
 sky130_fd_sc_hd__o2111ai_2 _17728_ (.A1(_08513_),
    .A2(_08516_),
    .B1(_08588_),
    .C1(_08589_),
    .D1(_08519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08591_));
 sky130_fd_sc_hd__a32o_2 _17729_ (.A1(_08518_),
    .A2(_08479_),
    .A3(_08517_),
    .B1(_08588_),
    .B2(_08589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08592_));
 sky130_fd_sc_hd__nand2_2 _17730_ (.A(_08591_),
    .B(_08592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08593_));
 sky130_fd_sc_hd__nand2_2 _17731_ (.A(\a_l[9] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08594_));
 sky130_fd_sc_hd__o2bb2ai_2 _17732_ (.A1_N(_08515_),
    .A2_N(_08512_),
    .B1(_08510_),
    .B2(_08507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08595_));
 sky130_fd_sc_hd__o21ai_2 _17733_ (.A1(_08482_),
    .A2(_08485_),
    .B1(_08595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08596_));
 sky130_fd_sc_hd__o2111ai_2 _17734_ (.A1(_02589_),
    .A2(_07234_),
    .B1(_08486_),
    .C1(_08511_),
    .D1(_08517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08597_));
 sky130_fd_sc_hd__a22o_2 _17735_ (.A1(\a_l[9] ),
    .A2(\b_h[15] ),
    .B1(_08596_),
    .B2(_08597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08598_));
 sky130_fd_sc_hd__nand4_2 _17736_ (.A(_08596_),
    .B(_08597_),
    .C(\a_l[9] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08599_));
 sky130_fd_sc_hd__a21o_2 _17737_ (.A1(_08596_),
    .A2(_08597_),
    .B1(_08594_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08600_));
 sky130_fd_sc_hd__o211ai_2 _17738_ (.A1(_09275_),
    .A2(_09679_),
    .B1(_08596_),
    .C1(_08597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08601_));
 sky130_fd_sc_hd__nand3_2 _17739_ (.A(_08593_),
    .B(_08598_),
    .C(_08599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08602_));
 sky130_fd_sc_hd__nand4_2 _17740_ (.A(_08591_),
    .B(_08592_),
    .C(_08600_),
    .D(_08601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08603_));
 sky130_fd_sc_hd__nand3_2 _17741_ (.A(_08593_),
    .B(_08600_),
    .C(_08601_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_2 _17742_ (.A(_08592_),
    .B(_08598_),
    .C(_08599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08605_));
 sky130_fd_sc_hd__nand4_2 _17743_ (.A(_08591_),
    .B(_08592_),
    .C(_08598_),
    .D(_08599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08606_));
 sky130_fd_sc_hd__nand3_2 _17744_ (.A(_08548_),
    .B(_08604_),
    .C(_08606_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08607_));
 sky130_fd_sc_hd__nand3_2 _17745_ (.A(_08549_),
    .B(_08602_),
    .C(_08603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08608_));
 sky130_fd_sc_hd__a22o_2 _17746_ (.A1(_08471_),
    .A2(_08473_),
    .B1(_08607_),
    .B2(_08608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08609_));
 sky130_fd_sc_hd__nand4_2 _17747_ (.A(_08471_),
    .B(_08473_),
    .C(_08607_),
    .D(_08608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08610_));
 sky130_fd_sc_hd__a21bo_2 _17748_ (.A1(_08533_),
    .A2(_08535_),
    .B1_N(_08534_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08611_));
 sky130_fd_sc_hd__a21oi_2 _17749_ (.A1(_08609_),
    .A2(_08610_),
    .B1(_08611_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08612_));
 sky130_fd_sc_hd__nand3_2 _17750_ (.A(_08611_),
    .B(_08610_),
    .C(_08609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08613_));
 sky130_fd_sc_hd__and2b_2 _17751_ (.A_N(_08612_),
    .B(_08613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08614_));
 sky130_fd_sc_hd__nand4_2 _17752_ (.A(_08456_),
    .B(_08457_),
    .C(_08541_),
    .D(_08542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08615_));
 sky130_fd_sc_hd__nand4_2 _17753_ (.A(_08543_),
    .B(_08460_),
    .C(_08457_),
    .D(_08456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08616_));
 sky130_fd_sc_hd__a21boi_2 _17754_ (.A1(_08457_),
    .A2(_08542_),
    .B1_N(_08541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08617_));
 sky130_fd_sc_hd__inv_2 _17755_ (.A(_08617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08618_));
 sky130_fd_sc_hd__o21bai_2 _17756_ (.A1(_08615_),
    .A2(_08459_),
    .B1_N(_08617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08619_));
 sky130_fd_sc_hd__nor3_2 _17757_ (.A(_08271_),
    .B(_08368_),
    .C(_08615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08620_));
 sky130_fd_sc_hd__nor2_2 _17758_ (.A(_08619_),
    .B(_08620_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08621_));
 sky130_fd_sc_hd__a21oi_2 _17759_ (.A1(_08274_),
    .A2(_08027_),
    .B1(_08619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08622_));
 sky130_fd_sc_hd__nand4_2 _17760_ (.A(_08278_),
    .B(_08616_),
    .C(_08618_),
    .D(_08273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08623_));
 sky130_fd_sc_hd__a21oi_2 _17761_ (.A1(_07587_),
    .A2(_08276_),
    .B1(_08623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08624_));
 sky130_fd_sc_hd__nand3_2 _17762_ (.A(_08277_),
    .B(_08622_),
    .C(_08273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08625_));
 sky130_fd_sc_hd__o21a_2 _17763_ (.A1(_08619_),
    .A2(_08620_),
    .B1(_08625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08626_));
 sky130_fd_sc_hd__o21ai_2 _17764_ (.A1(_08614_),
    .A2(_08626_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08627_));
 sky130_fd_sc_hd__a21oi_2 _17765_ (.A1(_08614_),
    .A2(_08626_),
    .B1(_08627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00362_));
 sky130_fd_sc_hd__and2_2 _17766_ (.A(_08596_),
    .B(_08599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08628_));
 sky130_fd_sc_hd__nand2_2 _17767_ (.A(\a_l[13] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08629_));
 sky130_fd_sc_hd__nand4_2 _17768_ (.A(\a_l[12] ),
    .B(\a_l[13] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08630_));
 sky130_fd_sc_hd__a22o_2 _17769_ (.A1(\a_l[13] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08631_));
 sky130_fd_sc_hd__a22o_2 _17770_ (.A1(\a_l[11] ),
    .A2(\b_h[14] ),
    .B1(_08630_),
    .B2(_08631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08632_));
 sky130_fd_sc_hd__nand4_2 _17771_ (.A(_08631_),
    .B(\b_h[14] ),
    .C(\a_l[11] ),
    .D(_08630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08633_));
 sky130_fd_sc_hd__o21ai_2 _17772_ (.A1(_08563_),
    .A2(_08566_),
    .B1(_08564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_2 _17773_ (.A(\a_l[15] ),
    .B(\b_h[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08635_));
 sky130_fd_sc_hd__a22o_2 _17774_ (.A1(\a_l[15] ),
    .A2(\b_h[10] ),
    .B1(\b_h[11] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08636_));
 sky130_fd_sc_hd__o21ai_2 _17775_ (.A1(_08494_),
    .A2(_08635_),
    .B1(_08636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08637_));
 sky130_fd_sc_hd__o211ai_2 _17776_ (.A1(_08566_),
    .A2(_08563_),
    .B1(_08564_),
    .C1(_08637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08638_));
 sky130_fd_sc_hd__o211a_2 _17777_ (.A1(_08494_),
    .A2(_08635_),
    .B1(_08636_),
    .C1(_08634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08639_));
 sky130_fd_sc_hd__o211ai_2 _17778_ (.A1(_08494_),
    .A2(_08635_),
    .B1(_08636_),
    .C1(_08634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08640_));
 sky130_fd_sc_hd__a22o_2 _17779_ (.A1(_08632_),
    .A2(_08633_),
    .B1(_08638_),
    .B2(_08640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08641_));
 sky130_fd_sc_hd__nand4_2 _17780_ (.A(_08632_),
    .B(_08633_),
    .C(_08638_),
    .D(_08640_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08642_));
 sky130_fd_sc_hd__nand2_2 _17781_ (.A(_08641_),
    .B(_08642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08643_));
 sky130_fd_sc_hd__o21ai_2 _17782_ (.A1(_08562_),
    .A2(_08574_),
    .B1(_08576_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08644_));
 sky130_fd_sc_hd__nand3_2 _17783_ (.A(_08644_),
    .B(_08642_),
    .C(_08641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08645_));
 sky130_fd_sc_hd__xnor2_2 _17784_ (.A(_08643_),
    .B(_08644_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08646_));
 sky130_fd_sc_hd__nand2_2 _17785_ (.A(\a_l[10] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08647_));
 sky130_fd_sc_hd__o31a_2 _17786_ (.A1(_09297_),
    .A2(_09657_),
    .A3(_08553_),
    .B1(_08558_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08648_));
 sky130_fd_sc_hd__o21bai_2 _17787_ (.A1(_08577_),
    .A2(_08585_),
    .B1_N(_08587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08649_));
 sky130_fd_sc_hd__o21ai_2 _17788_ (.A1(_08580_),
    .A2(_08583_),
    .B1(_08587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08650_));
 sky130_fd_sc_hd__and3_2 _17789_ (.A(_08586_),
    .B(_08650_),
    .C(_08648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08651_));
 sky130_fd_sc_hd__nand3_2 _17790_ (.A(_08586_),
    .B(_08650_),
    .C(_08648_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08652_));
 sky130_fd_sc_hd__o221ai_2 _17791_ (.A1(_08554_),
    .A2(_08557_),
    .B1(_08580_),
    .B2(_08583_),
    .C1(_08649_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08653_));
 sky130_fd_sc_hd__nand2_2 _17792_ (.A(_08652_),
    .B(_08653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08654_));
 sky130_fd_sc_hd__nand4_2 _17793_ (.A(_08652_),
    .B(_08653_),
    .C(\a_l[10] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08655_));
 sky130_fd_sc_hd__a22o_2 _17794_ (.A1(\a_l[10] ),
    .A2(\b_h[15] ),
    .B1(_08652_),
    .B2(_08653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08656_));
 sky130_fd_sc_hd__a21o_2 _17795_ (.A1(_08655_),
    .A2(_08656_),
    .B1(_08646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08657_));
 sky130_fd_sc_hd__a21boi_2 _17796_ (.A1(_08647_),
    .A2(_08654_),
    .B1_N(_08646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08658_));
 sky130_fd_sc_hd__nand3_2 _17797_ (.A(_08656_),
    .B(_08646_),
    .C(_08655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08659_));
 sky130_fd_sc_hd__nand2_2 _17798_ (.A(_08657_),
    .B(_08659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08660_));
 sky130_fd_sc_hd__o21ai_2 _17799_ (.A1(_08520_),
    .A2(_08590_),
    .B1(_08605_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08661_));
 sky130_fd_sc_hd__o211ai_2 _17800_ (.A1(_08520_),
    .A2(_08590_),
    .B1(_08605_),
    .C1(_08660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08662_));
 sky130_fd_sc_hd__nand3_2 _17801_ (.A(_08661_),
    .B(_08659_),
    .C(_08657_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08663_));
 sky130_fd_sc_hd__a21bo_2 _17802_ (.A1(_08662_),
    .A2(_08663_),
    .B1_N(_08628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08664_));
 sky130_fd_sc_hd__nand3b_2 _17803_ (.A_N(_08628_),
    .B(_08662_),
    .C(_08663_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08665_));
 sky130_fd_sc_hd__nand2_2 _17804_ (.A(_08607_),
    .B(_08610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08666_));
 sky130_fd_sc_hd__a21oi_2 _17805_ (.A1(_08664_),
    .A2(_08665_),
    .B1(_08666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08667_));
 sky130_fd_sc_hd__nand3_2 _17806_ (.A(_08666_),
    .B(_08665_),
    .C(_08664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08668_));
 sky130_fd_sc_hd__and2b_2 _17807_ (.A_N(_08667_),
    .B(_08668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08669_));
 sky130_fd_sc_hd__o31ai_2 _17808_ (.A1(_08612_),
    .A2(_08621_),
    .A3(_08624_),
    .B1(_08613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08670_));
 sky130_fd_sc_hd__a21oi_2 _17809_ (.A1(_08670_),
    .A2(_08669_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08671_));
 sky130_fd_sc_hd__o21a_2 _17810_ (.A1(_08669_),
    .A2(_08670_),
    .B1(_08671_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00363_));
 sky130_fd_sc_hd__a31oi_2 _17811_ (.A1(_08632_),
    .A2(_08633_),
    .A3(_08638_),
    .B1(_08639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08672_));
 sky130_fd_sc_hd__a21o_2 _17812_ (.A1(\a_l[14] ),
    .A2(\b_h[10] ),
    .B1(_09373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08673_));
 sky130_fd_sc_hd__and3_2 _17813_ (.A(_08494_),
    .B(\b_h[11] ),
    .C(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08674_));
 sky130_fd_sc_hd__and2_2 _17814_ (.A(\a_l[12] ),
    .B(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08675_));
 sky130_fd_sc_hd__nand2_2 _17815_ (.A(\a_l[14] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08676_));
 sky130_fd_sc_hd__nand2_2 _17816_ (.A(\a_l[13] ),
    .B(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08677_));
 sky130_fd_sc_hd__nand2_2 _17817_ (.A(\a_l[14] ),
    .B(\b_h[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08678_));
 sky130_fd_sc_hd__nand4_2 _17818_ (.A(\a_l[13] ),
    .B(\a_l[14] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08679_));
 sky130_fd_sc_hd__nand2_2 _17819_ (.A(_08677_),
    .B(_08678_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08680_));
 sky130_fd_sc_hd__and3_2 _17820_ (.A(_08680_),
    .B(_08675_),
    .C(_08679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08681_));
 sky130_fd_sc_hd__o2111ai_2 _17821_ (.A1(_08629_),
    .A2(_08676_),
    .B1(\a_l[12] ),
    .C1(\b_h[14] ),
    .D1(_08680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08682_));
 sky130_fd_sc_hd__a21oi_2 _17822_ (.A1(_08679_),
    .A2(_08680_),
    .B1(_08675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08683_));
 sky130_fd_sc_hd__o22ai_2 _17823_ (.A1(_09646_),
    .A2(_08673_),
    .B1(_08681_),
    .B2(_08683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08684_));
 sky130_fd_sc_hd__nand3b_2 _17824_ (.A_N(_08683_),
    .B(_08674_),
    .C(_08682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08685_));
 sky130_fd_sc_hd__nand2_2 _17825_ (.A(_08684_),
    .B(_08685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08686_));
 sky130_fd_sc_hd__xnor2_2 _17826_ (.A(_08672_),
    .B(_08686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08687_));
 sky130_fd_sc_hd__nand2_2 _17827_ (.A(\a_l[11] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08688_));
 sky130_fd_sc_hd__o31a_2 _17828_ (.A1(_09340_),
    .A2(_09657_),
    .A3(_08553_),
    .B1(_08633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08689_));
 sky130_fd_sc_hd__o21ai_2 _17829_ (.A1(_08553_),
    .A2(_08629_),
    .B1(_08633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_2 _17830_ (.A(_08645_),
    .B(_08689_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08691_));
 sky130_fd_sc_hd__inv_2 _17831_ (.A(_08691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08692_));
 sky130_fd_sc_hd__nand4_2 _17832_ (.A(_08644_),
    .B(_08690_),
    .C(_08641_),
    .D(_08642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08693_));
 sky130_fd_sc_hd__a22o_2 _17833_ (.A1(\a_l[11] ),
    .A2(\b_h[15] ),
    .B1(_08691_),
    .B2(_08693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08694_));
 sky130_fd_sc_hd__o21ai_2 _17834_ (.A1(_09297_),
    .A2(_09679_),
    .B1(_08693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08695_));
 sky130_fd_sc_hd__a21o_2 _17835_ (.A1(_08691_),
    .A2(_08693_),
    .B1(_08688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08696_));
 sky130_fd_sc_hd__o211ai_2 _17836_ (.A1(_08695_),
    .A2(_08692_),
    .B1(_08687_),
    .C1(_08696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08697_));
 sky130_fd_sc_hd__a41oi_2 _17837_ (.A1(\a_l[11] ),
    .A2(\b_h[15] ),
    .A3(_08691_),
    .A4(_08693_),
    .B1(_08687_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08698_));
 sky130_fd_sc_hd__nand2_2 _17838_ (.A(_08698_),
    .B(_08694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08699_));
 sky130_fd_sc_hd__nand2_2 _17839_ (.A(_08697_),
    .B(_08699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08700_));
 sky130_fd_sc_hd__nand4_2 _17840_ (.A(_08658_),
    .B(_08697_),
    .C(_08699_),
    .D(_08655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08701_));
 sky130_fd_sc_hd__nand2_2 _17841_ (.A(_08659_),
    .B(_08700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08702_));
 sky130_fd_sc_hd__o31a_2 _17842_ (.A1(_09286_),
    .A2(_09679_),
    .A3(_08651_),
    .B1(_08653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08703_));
 sky130_fd_sc_hd__a21o_2 _17843_ (.A1(_08701_),
    .A2(_08702_),
    .B1(_08703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08704_));
 sky130_fd_sc_hd__o2111ai_2 _17844_ (.A1(_08647_),
    .A2(_08651_),
    .B1(_08653_),
    .C1(_08701_),
    .D1(_08702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08705_));
 sky130_fd_sc_hd__nand2_2 _17845_ (.A(_08704_),
    .B(_08705_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08706_));
 sky130_fd_sc_hd__nand2_2 _17846_ (.A(_08663_),
    .B(_08628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08707_));
 sky130_fd_sc_hd__nand3_2 _17847_ (.A(_08706_),
    .B(_08707_),
    .C(_08662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08708_));
 sky130_fd_sc_hd__inv_2 _17848_ (.A(_08708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08709_));
 sky130_fd_sc_hd__a21o_2 _17849_ (.A1(_08662_),
    .A2(_08707_),
    .B1(_08706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08710_));
 sky130_fd_sc_hd__nand2_2 _17850_ (.A(_08708_),
    .B(_08710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08711_));
 sky130_fd_sc_hd__inv_2 _17851_ (.A(_08711_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08712_));
 sky130_fd_sc_hd__o211ai_2 _17852_ (.A1(_08619_),
    .A2(_08620_),
    .B1(_08669_),
    .C1(_08614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08713_));
 sky130_fd_sc_hd__a21oi_2 _17853_ (.A1(_08613_),
    .A2(_08668_),
    .B1(_08667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08714_));
 sky130_fd_sc_hd__o21bai_2 _17854_ (.A1(_08713_),
    .A2(_08624_),
    .B1_N(_08714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08715_));
 sky130_fd_sc_hd__nand2_2 _17855_ (.A(_08715_),
    .B(_08712_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08716_));
 sky130_fd_sc_hd__a21oi_2 _17856_ (.A1(_08715_),
    .A2(_08712_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08717_));
 sky130_fd_sc_hd__o21a_2 _17857_ (.A1(_08712_),
    .A2(_08715_),
    .B1(_08717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00364_));
 sky130_fd_sc_hd__nand4_2 _17858_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[12] ),
    .D(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08718_));
 sky130_fd_sc_hd__a22o_2 _17859_ (.A1(\a_l[15] ),
    .A2(\b_h[12] ),
    .B1(\b_h[13] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08719_));
 sky130_fd_sc_hd__and4_2 _17860_ (.A(_08719_),
    .B(\b_h[14] ),
    .C(\a_l[13] ),
    .D(_08718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08720_));
 sky130_fd_sc_hd__o2bb2a_2 _17861_ (.A1_N(_08718_),
    .A2_N(_08719_),
    .B1(_09340_),
    .B2(_09668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08721_));
 sky130_fd_sc_hd__nor2_2 _17862_ (.A(_08720_),
    .B(_08721_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08722_));
 sky130_fd_sc_hd__o21ai_2 _17863_ (.A1(_08494_),
    .A2(_08635_),
    .B1(_08685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08723_));
 sky130_fd_sc_hd__xnor2_2 _17864_ (.A(_08722_),
    .B(_08723_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08724_));
 sky130_fd_sc_hd__a41o_2 _17865_ (.A1(\a_l[13] ),
    .A2(\a_l[14] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_08681_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08725_));
 sky130_fd_sc_hd__o221ai_2 _17866_ (.A1(_08629_),
    .A2(_08676_),
    .B1(_08686_),
    .B2(_08672_),
    .C1(_08682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08726_));
 sky130_fd_sc_hd__nand4b_2 _17867_ (.A_N(_08672_),
    .B(_08684_),
    .C(_08685_),
    .D(_08725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08727_));
 sky130_fd_sc_hd__nand2_2 _17868_ (.A(_08726_),
    .B(_08727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08728_));
 sky130_fd_sc_hd__nand2_2 _17869_ (.A(\a_l[12] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08729_));
 sky130_fd_sc_hd__o2bb2a_2 _17870_ (.A1_N(_08726_),
    .A2_N(_08727_),
    .B1(_09319_),
    .B2(_09679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08730_));
 sky130_fd_sc_hd__and4_2 _17871_ (.A(_08726_),
    .B(_08727_),
    .C(\a_l[12] ),
    .D(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08731_));
 sky130_fd_sc_hd__o21ai_2 _17872_ (.A1(_08730_),
    .A2(_08731_),
    .B1(_08724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08732_));
 sky130_fd_sc_hd__a21oi_2 _17873_ (.A1(_08728_),
    .A2(_08729_),
    .B1(_08724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08733_));
 sky130_fd_sc_hd__o21ai_2 _17874_ (.A1(_08728_),
    .A2(_08729_),
    .B1(_08733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08734_));
 sky130_fd_sc_hd__nand2_2 _17875_ (.A(_08732_),
    .B(_08734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08735_));
 sky130_fd_sc_hd__a22oi_2 _17876_ (.A1(_08694_),
    .A2(_08698_),
    .B1(_08732_),
    .B2(_08734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08736_));
 sky130_fd_sc_hd__and4_2 _17877_ (.A(_08694_),
    .B(_08732_),
    .C(_08734_),
    .D(_08698_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08737_));
 sky130_fd_sc_hd__o31a_2 _17878_ (.A1(_09297_),
    .A2(_09679_),
    .A3(_08692_),
    .B1(_08693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08738_));
 sky130_fd_sc_hd__o21ai_2 _17879_ (.A1(_08736_),
    .A2(_08737_),
    .B1(_08738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08739_));
 sky130_fd_sc_hd__a21o_2 _17880_ (.A1(_08699_),
    .A2(_08735_),
    .B1(_08738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08740_));
 sky130_fd_sc_hd__o21ai_2 _17881_ (.A1(_08737_),
    .A2(_08740_),
    .B1(_08739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08741_));
 sky130_fd_sc_hd__a21boi_2 _17882_ (.A1(_08701_),
    .A2(_08703_),
    .B1_N(_08702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08742_));
 sky130_fd_sc_hd__nand2b_2 _17883_ (.A_N(_08742_),
    .B(_08741_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08743_));
 sky130_fd_sc_hd__o211a_2 _17884_ (.A1(_08737_),
    .A2(_08740_),
    .B1(_08742_),
    .C1(_08739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08744_));
 sky130_fd_sc_hd__o211ai_2 _17885_ (.A1(_08737_),
    .A2(_08740_),
    .B1(_08742_),
    .C1(_08739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08745_));
 sky130_fd_sc_hd__nand2_2 _17886_ (.A(_08743_),
    .B(_08745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08746_));
 sky130_fd_sc_hd__inv_2 _17887_ (.A(_08746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08747_));
 sky130_fd_sc_hd__a211oi_2 _17888_ (.A1(_08715_),
    .A2(_08712_),
    .B1(_08709_),
    .C1(_08747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08748_));
 sky130_fd_sc_hd__a21oi_2 _17889_ (.A1(_08708_),
    .A2(_08716_),
    .B1(_08746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08749_));
 sky130_fd_sc_hd__nor3_2 _17890_ (.A(rst),
    .B(_08748_),
    .C(_08749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00365_));
 sky130_fd_sc_hd__a41o_2 _17891_ (.A1(\a_l[14] ),
    .A2(\a_l[15] ),
    .A3(\b_h[12] ),
    .A4(\b_h[13] ),
    .B1(_08720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08750_));
 sky130_fd_sc_hd__a21oi_2 _17892_ (.A1(_08723_),
    .A2(_08722_),
    .B1(_08750_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08751_));
 sky130_fd_sc_hd__and3_2 _17893_ (.A(_08723_),
    .B(_08750_),
    .C(_08722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08752_));
 sky130_fd_sc_hd__nor4_2 _17894_ (.A(_09340_),
    .B(_09679_),
    .C(_08751_),
    .D(_08752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08753_));
 sky130_fd_sc_hd__o22a_2 _17895_ (.A1(_09340_),
    .A2(_09679_),
    .B1(_08751_),
    .B2(_08752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08754_));
 sky130_fd_sc_hd__a22o_2 _17896_ (.A1(\a_l[15] ),
    .A2(\b_h[13] ),
    .B1(\b_h[14] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08755_));
 sky130_fd_sc_hd__nand4_2 _17897_ (.A(\a_l[14] ),
    .B(\a_l[15] ),
    .C(\b_h[13] ),
    .D(\b_h[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_2 _17898_ (.A(_08755_),
    .B(_08756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08757_));
 sky130_fd_sc_hd__and4bb_2 _17899_ (.A_N(_08753_),
    .B_N(_08754_),
    .C(_08755_),
    .D(_08756_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08758_));
 sky130_fd_sc_hd__o21a_2 _17900_ (.A1(_08753_),
    .A2(_08754_),
    .B1(_08757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08759_));
 sky130_fd_sc_hd__nor2_2 _17901_ (.A(_08758_),
    .B(_08759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08760_));
 sky130_fd_sc_hd__o311a_2 _17902_ (.A1(_09319_),
    .A2(_09679_),
    .A3(_08728_),
    .B1(_08733_),
    .C1(_08760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08761_));
 sky130_fd_sc_hd__xor2_2 _17903_ (.A(_08734_),
    .B(_08760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08762_));
 sky130_fd_sc_hd__or3b_2 _17904_ (.A(_09319_),
    .B(_09679_),
    .C_N(_08726_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08763_));
 sky130_fd_sc_hd__and2_2 _17905_ (.A(_08762_),
    .B(_08763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08764_));
 sky130_fd_sc_hd__a21oi_2 _17906_ (.A1(_08727_),
    .A2(_08763_),
    .B1(_08762_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08765_));
 sky130_fd_sc_hd__a21o_2 _17907_ (.A1(_08764_),
    .A2(_08727_),
    .B1(_08765_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08766_));
 sky130_fd_sc_hd__o21ai_2 _17908_ (.A1(_08699_),
    .A2(_08735_),
    .B1(_08740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08767_));
 sky130_fd_sc_hd__inv_2 _17909_ (.A(_08767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08768_));
 sky130_fd_sc_hd__nor2_2 _17910_ (.A(_08768_),
    .B(_08766_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08769_));
 sky130_fd_sc_hd__xnor2_2 _17911_ (.A(_08766_),
    .B(_08768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08770_));
 sky130_fd_sc_hd__nor2_2 _17912_ (.A(_08711_),
    .B(_08746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08771_));
 sky130_fd_sc_hd__and3_2 _17913_ (.A(_08614_),
    .B(_08669_),
    .C(_08771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08772_));
 sky130_fd_sc_hd__o21a_2 _17914_ (.A1(_08619_),
    .A2(_08620_),
    .B1(_08772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08773_));
 sky130_fd_sc_hd__o21ai_2 _17915_ (.A1(_08619_),
    .A2(_08620_),
    .B1(_08772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08774_));
 sky130_fd_sc_hd__a221o_2 _17916_ (.A1(_08709_),
    .A2(_08743_),
    .B1(_08771_),
    .B2(_08714_),
    .C1(_08744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08775_));
 sky130_fd_sc_hd__o21bai_2 _17917_ (.A1(_08774_),
    .A2(_08624_),
    .B1_N(_08775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08776_));
 sky130_fd_sc_hd__a21oi_2 _17918_ (.A1(_08625_),
    .A2(_08773_),
    .B1(_08775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08777_));
 sky130_fd_sc_hd__o21ai_2 _17919_ (.A1(_08770_),
    .A2(_08777_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08778_));
 sky130_fd_sc_hd__a21oi_2 _17920_ (.A1(_08770_),
    .A2(_08777_),
    .B1(_08778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00366_));
 sky130_fd_sc_hd__a31o_2 _17921_ (.A1(_08722_),
    .A2(_08723_),
    .A3(_08750_),
    .B1(_08753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08779_));
 sky130_fd_sc_hd__nand2_2 _17922_ (.A(\a_l[14] ),
    .B(\b_h[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08780_));
 sky130_fd_sc_hd__o22a_2 _17923_ (.A1(\b_h[15] ),
    .A2(_08676_),
    .B1(_08780_),
    .B2(\b_h[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08781_));
 sky130_fd_sc_hd__or3_2 _17924_ (.A(_09373_),
    .B(_09668_),
    .C(_08781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08782_));
 sky130_fd_sc_hd__a22o_2 _17925_ (.A1(\a_l[15] ),
    .A2(\b_h[14] ),
    .B1(\b_h[15] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08783_));
 sky130_fd_sc_hd__a21oi_2 _17926_ (.A1(_08782_),
    .A2(_08783_),
    .B1(_08758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08784_));
 sky130_fd_sc_hd__o311a_2 _17927_ (.A1(_09373_),
    .A2(_09668_),
    .A3(_08781_),
    .B1(_08783_),
    .C1(_08758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08785_));
 sky130_fd_sc_hd__nor2_2 _17928_ (.A(_08784_),
    .B(_08785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08786_));
 sky130_fd_sc_hd__xnor2_2 _17929_ (.A(_08779_),
    .B(_08786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08787_));
 sky130_fd_sc_hd__o21ba_2 _17930_ (.A1(_08761_),
    .A2(_08765_),
    .B1_N(_08787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08788_));
 sky130_fd_sc_hd__or3b_2 _17931_ (.A(_08761_),
    .B(_08765_),
    .C_N(_08787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08789_));
 sky130_fd_sc_hd__inv_2 _17932_ (.A(_08789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08790_));
 sky130_fd_sc_hd__nand2b_2 _17933_ (.A_N(_08788_),
    .B(_08789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08791_));
 sky130_fd_sc_hd__inv_2 _17934_ (.A(_08791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08792_));
 sky130_fd_sc_hd__o22ai_2 _17935_ (.A1(_08766_),
    .A2(_08768_),
    .B1(_08770_),
    .B2(_08777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08793_));
 sky130_fd_sc_hd__o22ai_2 _17936_ (.A1(_08788_),
    .A2(_08790_),
    .B1(_08770_),
    .B2(_08777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_2 _17937_ (.A(_08793_),
    .B(_08792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08795_));
 sky130_fd_sc_hd__o211a_2 _17938_ (.A1(_08794_),
    .A2(_08769_),
    .B1(_09690_),
    .C1(_08795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00367_));
 sky130_fd_sc_hd__o21a_2 _17939_ (.A1(_09373_),
    .A2(_09679_),
    .B1(_08782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08796_));
 sky130_fd_sc_hd__a41o_2 _17940_ (.A1(\a_l[14] ),
    .A2(\a_l[15] ),
    .A3(\b_h[14] ),
    .A4(\b_h[15] ),
    .B1(_08796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08797_));
 sky130_fd_sc_hd__a21oi_2 _17941_ (.A1(_08786_),
    .A2(_08779_),
    .B1(_08785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08798_));
 sky130_fd_sc_hd__xor2_2 _17942_ (.A(_08797_),
    .B(_08798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08799_));
 sky130_fd_sc_hd__inv_2 _17943_ (.A(_08799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08800_));
 sky130_fd_sc_hd__nor2_2 _17944_ (.A(_08769_),
    .B(_08788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08801_));
 sky130_fd_sc_hd__o21a_2 _17945_ (.A1(_08769_),
    .A2(_08788_),
    .B1(_08789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08802_));
 sky130_fd_sc_hd__o21ai_2 _17946_ (.A1(_08769_),
    .A2(_08788_),
    .B1(_08789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08803_));
 sky130_fd_sc_hd__nor2_2 _17947_ (.A(_08770_),
    .B(_08791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08804_));
 sky130_fd_sc_hd__or2_2 _17948_ (.A(_08770_),
    .B(_08791_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08805_));
 sky130_fd_sc_hd__nand2_2 _17949_ (.A(_08776_),
    .B(_08804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08806_));
 sky130_fd_sc_hd__o22ai_2 _17950_ (.A1(_08790_),
    .A2(_08801_),
    .B1(_08805_),
    .B2(_08777_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08807_));
 sky130_fd_sc_hd__a211oi_2 _17951_ (.A1(_08776_),
    .A2(_08804_),
    .B1(_08802_),
    .C1(_08799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08808_));
 sky130_fd_sc_hd__a21oi_2 _17952_ (.A1(_08803_),
    .A2(_08806_),
    .B1(_08800_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08809_));
 sky130_fd_sc_hd__nand2_2 _17953_ (.A(_08807_),
    .B(_08799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08810_));
 sky130_fd_sc_hd__nor3_2 _17954_ (.A(rst),
    .B(_08808_),
    .C(_08809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00368_));
 sky130_fd_sc_hd__o32a_2 _17955_ (.A1(_09373_),
    .A2(_09668_),
    .A3(_08780_),
    .B1(_08796_),
    .B2(_08798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08811_));
 sky130_fd_sc_hd__a21oi_2 _17956_ (.A1(_08810_),
    .A2(_08811_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00369_));
 sky130_fd_sc_hd__and3_2 _17957_ (.A(_09690_),
    .B(\a_l[0] ),
    .C(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00370_));
 sky130_fd_sc_hd__a22oi_2 _17958_ (.A1(\b_l[0] ),
    .A2(\a_l[1] ),
    .B1(\a_l[0] ),
    .B2(\b_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08812_));
 sky130_fd_sc_hd__a311oi_2 _17959_ (.A1(\a_l[1] ),
    .A2(\a_l[0] ),
    .A3(_04133_),
    .B1(_08812_),
    .C1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00371_));
 sky130_fd_sc_hd__and3_2 _17960_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(_04133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08813_));
 sky130_fd_sc_hd__a22oi_2 _17961_ (.A1(\a_l[2] ),
    .A2(\b_l[0] ),
    .B1(\b_l[1] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08814_));
 sky130_fd_sc_hd__a211o_2 _17962_ (.A1(\b_l[2] ),
    .A2(\a_l[0] ),
    .B1(_08813_),
    .C1(_08814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08815_));
 sky130_fd_sc_hd__o211ai_2 _17963_ (.A1(_08813_),
    .A2(_08814_),
    .B1(\b_l[2] ),
    .C1(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08816_));
 sky130_fd_sc_hd__o211a_2 _17964_ (.A1(_04134_),
    .A2(_06402_),
    .B1(_08815_),
    .C1(_08816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08817_));
 sky130_fd_sc_hd__a211oi_2 _17965_ (.A1(_08815_),
    .A2(_08816_),
    .B1(_04134_),
    .C1(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08818_));
 sky130_fd_sc_hd__nor3_2 _17966_ (.A(rst),
    .B(_08817_),
    .C(_08818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00372_));
 sky130_fd_sc_hd__a22o_2 _17967_ (.A1(\a_l[2] ),
    .A2(\b_l[1] ),
    .B1(\a_l[3] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08819_));
 sky130_fd_sc_hd__and4_2 _17968_ (.A(\a_l[2] ),
    .B(\b_l[0] ),
    .C(\b_l[1] ),
    .D(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08820_));
 sky130_fd_sc_hd__nand4_2 _17969_ (.A(\a_l[2] ),
    .B(\b_l[0] ),
    .C(\b_l[1] ),
    .D(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08821_));
 sky130_fd_sc_hd__a22o_2 _17970_ (.A1(\a_l[1] ),
    .A2(\b_l[2] ),
    .B1(_08819_),
    .B2(_08821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08822_));
 sky130_fd_sc_hd__nand4_2 _17971_ (.A(_08819_),
    .B(_08821_),
    .C(\a_l[1] ),
    .D(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08823_));
 sky130_fd_sc_hd__o32ai_2 _17972_ (.A1(_09155_),
    .A2(_09166_),
    .A3(_08814_),
    .B1(_06441_),
    .B2(_04134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08824_));
 sky130_fd_sc_hd__a21o_2 _17973_ (.A1(_08822_),
    .A2(_08823_),
    .B1(_08824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08825_));
 sky130_fd_sc_hd__nand3_2 _17974_ (.A(_08824_),
    .B(_08823_),
    .C(_08822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08826_));
 sky130_fd_sc_hd__a22oi_2 _17975_ (.A1(\a_l[0] ),
    .A2(\b_l[3] ),
    .B1(_08825_),
    .B2(_08826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08827_));
 sky130_fd_sc_hd__and4_2 _17976_ (.A(_08825_),
    .B(_08826_),
    .C(\a_l[0] ),
    .D(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08828_));
 sky130_fd_sc_hd__nor2_2 _17977_ (.A(_08827_),
    .B(_08828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08829_));
 sky130_fd_sc_hd__a21oi_2 _17978_ (.A1(_08818_),
    .A2(_08829_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08830_));
 sky130_fd_sc_hd__o21a_2 _17979_ (.A1(_08818_),
    .A2(_08829_),
    .B1(_08830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00373_));
 sky130_fd_sc_hd__and3_2 _17980_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08831_));
 sky130_fd_sc_hd__a22oi_2 _17981_ (.A1(\a_l[1] ),
    .A2(\b_l[3] ),
    .B1(\b_l[4] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08832_));
 sky130_fd_sc_hd__nor2_2 _17982_ (.A(_08831_),
    .B(_08832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08833_));
 sky130_fd_sc_hd__a31o_2 _17983_ (.A1(\b_l[3] ),
    .A2(\b_l[4] ),
    .A3(_06401_),
    .B1(_08832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08834_));
 sky130_fd_sc_hd__a31oi_2 _17984_ (.A1(_08819_),
    .A2(\b_l[2] ),
    .A3(\a_l[1] ),
    .B1(_08820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08835_));
 sky130_fd_sc_hd__a31o_2 _17985_ (.A1(_08819_),
    .A2(\b_l[2] ),
    .A3(\a_l[1] ),
    .B1(_08820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08836_));
 sky130_fd_sc_hd__nand2_2 _17986_ (.A(\a_l[2] ),
    .B(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08837_));
 sky130_fd_sc_hd__and4_2 _17987_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[3] ),
    .D(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08838_));
 sky130_fd_sc_hd__nand4_2 _17988_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[3] ),
    .D(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08839_));
 sky130_fd_sc_hd__a22oi_2 _17989_ (.A1(\b_l[1] ),
    .A2(\a_l[3] ),
    .B1(\a_l[4] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08840_));
 sky130_fd_sc_hd__a22o_2 _17990_ (.A1(\b_l[1] ),
    .A2(\a_l[3] ),
    .B1(\a_l[4] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08841_));
 sky130_fd_sc_hd__o221ai_2 _17991_ (.A1(_09144_),
    .A2(_09155_),
    .B1(_04134_),
    .B2(_06521_),
    .C1(_08841_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08842_));
 sky130_fd_sc_hd__a21o_2 _17992_ (.A1(_08839_),
    .A2(_08841_),
    .B1(_08837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08843_));
 sky130_fd_sc_hd__o22a_2 _17993_ (.A1(_09144_),
    .A2(_09155_),
    .B1(_08838_),
    .B2(_08840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08844_));
 sky130_fd_sc_hd__o31ai_2 _17994_ (.A1(_08837_),
    .A2(_08838_),
    .A3(_08840_),
    .B1(_08836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08845_));
 sky130_fd_sc_hd__nand3_2 _17995_ (.A(_08843_),
    .B(_08835_),
    .C(_08842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08846_));
 sky130_fd_sc_hd__o21ai_2 _17996_ (.A1(_08844_),
    .A2(_08845_),
    .B1(_08846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08847_));
 sky130_fd_sc_hd__nand2_2 _17997_ (.A(_08847_),
    .B(_08833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08848_));
 sky130_fd_sc_hd__or2_2 _17998_ (.A(_08833_),
    .B(_08847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08849_));
 sky130_fd_sc_hd__nand3_2 _17999_ (.A(_08825_),
    .B(\b_l[3] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08850_));
 sky130_fd_sc_hd__and4_2 _18000_ (.A(_08826_),
    .B(_08848_),
    .C(_08849_),
    .D(_08850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08851_));
 sky130_fd_sc_hd__a22oi_2 _18001_ (.A1(_08834_),
    .A2(_08847_),
    .B1(_08850_),
    .B2(_08826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08852_));
 sky130_fd_sc_hd__o21ai_2 _18002_ (.A1(_08834_),
    .A2(_08847_),
    .B1(_08852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08853_));
 sky130_fd_sc_hd__and2b_2 _18003_ (.A_N(_08851_),
    .B(_08853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08854_));
 sky130_fd_sc_hd__a21o_2 _18004_ (.A1(_08818_),
    .A2(_08829_),
    .B1(_08854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08855_));
 sky130_fd_sc_hd__nand4b_2 _18005_ (.A_N(_08851_),
    .B(_08853_),
    .C(_08818_),
    .D(_08829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08856_));
 sky130_fd_sc_hd__and3_2 _18006_ (.A(_09690_),
    .B(_08855_),
    .C(_08856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00374_));
 sky130_fd_sc_hd__o2bb2ai_2 _18007_ (.A1_N(_08833_),
    .A2_N(_08846_),
    .B1(_08844_),
    .B2(_08845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08857_));
 sky130_fd_sc_hd__nand2_2 _18008_ (.A(\a_l[0] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08858_));
 sky130_fd_sc_hd__nand2_2 _18009_ (.A(\a_l[1] ),
    .B(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08859_));
 sky130_fd_sc_hd__nand2_2 _18010_ (.A(\a_l[2] ),
    .B(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08860_));
 sky130_fd_sc_hd__nand2_2 _18011_ (.A(_08859_),
    .B(_08860_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08861_));
 sky130_fd_sc_hd__o21ai_2 _18012_ (.A1(_04182_),
    .A2(_06441_),
    .B1(_08861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08862_));
 sky130_fd_sc_hd__o2111ai_2 _18013_ (.A1(_04182_),
    .A2(_06441_),
    .B1(\a_l[0] ),
    .C1(\b_l[5] ),
    .D1(_08861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08863_));
 sky130_fd_sc_hd__o21ai_2 _18014_ (.A1(_09166_),
    .A2(_09220_),
    .B1(_08862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08864_));
 sky130_fd_sc_hd__nand2_2 _18015_ (.A(_08863_),
    .B(_08864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08865_));
 sky130_fd_sc_hd__o21a_2 _18016_ (.A1(_04134_),
    .A2(_06521_),
    .B1(_08837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08866_));
 sky130_fd_sc_hd__o21ai_2 _18017_ (.A1(_08837_),
    .A2(_08840_),
    .B1(_08839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08867_));
 sky130_fd_sc_hd__o22a_2 _18018_ (.A1(_04134_),
    .A2(_06521_),
    .B1(_08837_),
    .B2(_08840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08868_));
 sky130_fd_sc_hd__nand2_2 _18019_ (.A(\b_l[2] ),
    .B(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08869_));
 sky130_fd_sc_hd__nand2_2 _18020_ (.A(\b_l[1] ),
    .B(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08870_));
 sky130_fd_sc_hd__nand2_2 _18021_ (.A(\b_l[0] ),
    .B(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08871_));
 sky130_fd_sc_hd__a22oi_2 _18022_ (.A1(\b_l[1] ),
    .A2(\a_l[4] ),
    .B1(\a_l[5] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08872_));
 sky130_fd_sc_hd__nand2_2 _18023_ (.A(_08870_),
    .B(_08871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08873_));
 sky130_fd_sc_hd__nand4_2 _18024_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[4] ),
    .D(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08874_));
 sky130_fd_sc_hd__nand4_2 _18025_ (.A(_08873_),
    .B(_08874_),
    .C(\b_l[2] ),
    .D(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08875_));
 sky130_fd_sc_hd__o2bb2ai_2 _18026_ (.A1_N(_08873_),
    .A2_N(_08874_),
    .B1(_09155_),
    .B2(_09188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08876_));
 sky130_fd_sc_hd__a21o_2 _18027_ (.A1(_08873_),
    .A2(_08874_),
    .B1(_08869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08877_));
 sky130_fd_sc_hd__o211ai_2 _18028_ (.A1(_09155_),
    .A2(_09188_),
    .B1(_08873_),
    .C1(_08874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08878_));
 sky130_fd_sc_hd__nand3_2 _18029_ (.A(_08876_),
    .B(_08867_),
    .C(_08875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08879_));
 sky130_fd_sc_hd__a2bb2oi_2 _18030_ (.A1_N(_08840_),
    .A2_N(_08866_),
    .B1(_08875_),
    .B2(_08876_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08880_));
 sky130_fd_sc_hd__nand3_2 _18031_ (.A(_08868_),
    .B(_08877_),
    .C(_08878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08881_));
 sky130_fd_sc_hd__a21o_2 _18032_ (.A1(_08879_),
    .A2(_08881_),
    .B1(_08865_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08882_));
 sky130_fd_sc_hd__nand3_2 _18033_ (.A(_08865_),
    .B(_08879_),
    .C(_08881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08883_));
 sky130_fd_sc_hd__nand2_2 _18034_ (.A(_08882_),
    .B(_08883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08884_));
 sky130_fd_sc_hd__a21boi_2 _18035_ (.A1(_08882_),
    .A2(_08883_),
    .B1_N(_08857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08885_));
 sky130_fd_sc_hd__nand2_2 _18036_ (.A(_08884_),
    .B(_08857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08886_));
 sky130_fd_sc_hd__nand3b_2 _18037_ (.A_N(_08857_),
    .B(_08882_),
    .C(_08883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08887_));
 sky130_fd_sc_hd__o2bb2ai_2 _18038_ (.A1_N(_08886_),
    .A2_N(_08887_),
    .B1(_04182_),
    .B2(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08888_));
 sky130_fd_sc_hd__nand3_2 _18039_ (.A(_08886_),
    .B(_08887_),
    .C(_08831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08889_));
 sky130_fd_sc_hd__nand2_2 _18040_ (.A(_08888_),
    .B(_08889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08890_));
 sky130_fd_sc_hd__nand3_2 _18041_ (.A(_08853_),
    .B(_08856_),
    .C(_08890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08891_));
 sky130_fd_sc_hd__nor2_2 _18042_ (.A(_08856_),
    .B(_08890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08892_));
 sky130_fd_sc_hd__nand3b_2 _18043_ (.A_N(_08853_),
    .B(_08888_),
    .C(_08889_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08893_));
 sky130_fd_sc_hd__a21o_2 _18044_ (.A1(_08853_),
    .A2(_08856_),
    .B1(_08890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08894_));
 sky130_fd_sc_hd__and3_2 _18045_ (.A(_09690_),
    .B(_08891_),
    .C(_08894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00375_));
 sky130_fd_sc_hd__nand2_2 _18046_ (.A(\a_l[0] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08895_));
 sky130_fd_sc_hd__o22a_2 _18047_ (.A1(_04182_),
    .A2(_06441_),
    .B1(_08858_),
    .B2(_08862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08896_));
 sky130_fd_sc_hd__o211a_2 _18048_ (.A1(_04182_),
    .A2(_06441_),
    .B1(_08863_),
    .C1(_08895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08897_));
 sky130_fd_sc_hd__nor2_2 _18049_ (.A(_08895_),
    .B(_08896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08898_));
 sky130_fd_sc_hd__nor2_2 _18050_ (.A(_08897_),
    .B(_08898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08899_));
 sky130_fd_sc_hd__inv_2 _18051_ (.A(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08900_));
 sky130_fd_sc_hd__a32oi_2 _18052_ (.A1(_08876_),
    .A2(_08867_),
    .A3(_08875_),
    .B1(_08864_),
    .B2(_08863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08901_));
 sky130_fd_sc_hd__a32o_2 _18053_ (.A1(_08876_),
    .A2(_08867_),
    .A3(_08875_),
    .B1(_08864_),
    .B2(_08863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08902_));
 sky130_fd_sc_hd__o21ai_2 _18054_ (.A1(_08865_),
    .A2(_08880_),
    .B1(_08879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08903_));
 sky130_fd_sc_hd__nand2_2 _18055_ (.A(\a_l[1] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08904_));
 sky130_fd_sc_hd__nand2_2 _18056_ (.A(\a_l[2] ),
    .B(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08905_));
 sky130_fd_sc_hd__nand2_2 _18057_ (.A(\a_l[3] ),
    .B(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08906_));
 sky130_fd_sc_hd__a22oi_2 _18058_ (.A1(\a_l[3] ),
    .A2(\b_l[3] ),
    .B1(\b_l[4] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_2 _18059_ (.A(_08905_),
    .B(_08906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08908_));
 sky130_fd_sc_hd__nand4_2 _18060_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_l[3] ),
    .D(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08909_));
 sky130_fd_sc_hd__a22oi_2 _18061_ (.A1(\a_l[1] ),
    .A2(\b_l[5] ),
    .B1(_08908_),
    .B2(_08909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08910_));
 sky130_fd_sc_hd__nand3_2 _18062_ (.A(_08909_),
    .B(\b_l[5] ),
    .C(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08911_));
 sky130_fd_sc_hd__a21oi_2 _18063_ (.A1(_08905_),
    .A2(_08906_),
    .B1(_08911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08912_));
 sky130_fd_sc_hd__nor2_2 _18064_ (.A(_08910_),
    .B(_08912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08913_));
 sky130_fd_sc_hd__o21ai_2 _18065_ (.A1(_08869_),
    .A2(_08872_),
    .B1(_08874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08914_));
 sky130_fd_sc_hd__o21a_2 _18066_ (.A1(_08869_),
    .A2(_08872_),
    .B1(_08874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08915_));
 sky130_fd_sc_hd__nand2_2 _18067_ (.A(\b_l[2] ),
    .B(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_2 _18068_ (.A(\b_l[0] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08917_));
 sky130_fd_sc_hd__nand2_2 _18069_ (.A(\b_l[1] ),
    .B(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08918_));
 sky130_fd_sc_hd__a22oi_2 _18070_ (.A1(\b_l[1] ),
    .A2(\a_l[5] ),
    .B1(\a_l[6] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08919_));
 sky130_fd_sc_hd__nand2_2 _18071_ (.A(_08917_),
    .B(_08918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08920_));
 sky130_fd_sc_hd__nand4_2 _18072_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[5] ),
    .D(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08921_));
 sky130_fd_sc_hd__and4_2 _18073_ (.A(_08920_),
    .B(_08921_),
    .C(\b_l[2] ),
    .D(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08922_));
 sky130_fd_sc_hd__o2111ai_2 _18074_ (.A1(_04134_),
    .A2(_06681_),
    .B1(\b_l[2] ),
    .C1(\a_l[4] ),
    .D1(_08920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08923_));
 sky130_fd_sc_hd__a22o_2 _18075_ (.A1(\b_l[2] ),
    .A2(\a_l[4] ),
    .B1(_08920_),
    .B2(_08921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08924_));
 sky130_fd_sc_hd__a21o_2 _18076_ (.A1(_08920_),
    .A2(_08921_),
    .B1(_08916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08925_));
 sky130_fd_sc_hd__o221ai_2 _18077_ (.A1(_09155_),
    .A2(_09199_),
    .B1(_04134_),
    .B2(_06681_),
    .C1(_08920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08926_));
 sky130_fd_sc_hd__nand2_2 _18078_ (.A(_08924_),
    .B(_08914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08927_));
 sky130_fd_sc_hd__nand3_2 _18079_ (.A(_08924_),
    .B(_08914_),
    .C(_08923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08928_));
 sky130_fd_sc_hd__nand3_2 _18080_ (.A(_08915_),
    .B(_08925_),
    .C(_08926_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08929_));
 sky130_fd_sc_hd__nand2_2 _18081_ (.A(_08928_),
    .B(_08929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08930_));
 sky130_fd_sc_hd__o211ai_2 _18082_ (.A1(_08910_),
    .A2(_08912_),
    .B1(_08928_),
    .C1(_08929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_2 _18083_ (.A(_08930_),
    .B(_08913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08932_));
 sky130_fd_sc_hd__a22oi_2 _18084_ (.A1(_08930_),
    .A2(_08913_),
    .B1(_08902_),
    .B2(_08881_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08933_));
 sky130_fd_sc_hd__o211a_2 _18085_ (.A1(_08880_),
    .A2(_08901_),
    .B1(_08931_),
    .C1(_08932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08934_));
 sky130_fd_sc_hd__o2111ai_2 _18086_ (.A1(_08880_),
    .A2(_08865_),
    .B1(_08879_),
    .C1(_08931_),
    .D1(_08932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08935_));
 sky130_fd_sc_hd__o21ai_2 _18087_ (.A1(_08910_),
    .A2(_08912_),
    .B1(_08930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08936_));
 sky130_fd_sc_hd__o211ai_2 _18088_ (.A1(_08922_),
    .A2(_08927_),
    .B1(_08929_),
    .C1(_08913_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08937_));
 sky130_fd_sc_hd__nand3_2 _18089_ (.A(_08936_),
    .B(_08937_),
    .C(_08903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08938_));
 sky130_fd_sc_hd__a21oi_2 _18090_ (.A1(_08935_),
    .A2(_08938_),
    .B1(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08939_));
 sky130_fd_sc_hd__a21o_2 _18091_ (.A1(_08935_),
    .A2(_08938_),
    .B1(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08940_));
 sky130_fd_sc_hd__and3_2 _18092_ (.A(_08935_),
    .B(_08938_),
    .C(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08941_));
 sky130_fd_sc_hd__nand3_2 _18093_ (.A(_08935_),
    .B(_08938_),
    .C(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08942_));
 sky130_fd_sc_hd__nand2_2 _18094_ (.A(_08940_),
    .B(_08942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08943_));
 sky130_fd_sc_hd__a21o_2 _18095_ (.A1(_08887_),
    .A2(_08831_),
    .B1(_08885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08944_));
 sky130_fd_sc_hd__a21oi_2 _18096_ (.A1(_08887_),
    .A2(_08831_),
    .B1(_08885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08945_));
 sky130_fd_sc_hd__a21oi_2 _18097_ (.A1(_08940_),
    .A2(_08942_),
    .B1(_08944_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08946_));
 sky130_fd_sc_hd__a221o_2 _18098_ (.A1(_08831_),
    .A2(_08887_),
    .B1(_08940_),
    .B2(_08942_),
    .C1(_08885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08947_));
 sky130_fd_sc_hd__nor3_2 _18099_ (.A(_08939_),
    .B(_08941_),
    .C(_08945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08948_));
 sky130_fd_sc_hd__or3_2 _18100_ (.A(_08939_),
    .B(_08941_),
    .C(_08945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08949_));
 sky130_fd_sc_hd__or2_2 _18101_ (.A(_08946_),
    .B(_08948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08950_));
 sky130_fd_sc_hd__nor3_2 _18102_ (.A(_08893_),
    .B(_08946_),
    .C(_08948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08951_));
 sky130_fd_sc_hd__o31a_2 _18103_ (.A1(_08946_),
    .A2(_08948_),
    .A3(_08894_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08952_));
 sky130_fd_sc_hd__a21boi_2 _18104_ (.A1(_08894_),
    .A2(_08950_),
    .B1_N(_08952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00376_));
 sky130_fd_sc_hd__a31oi_2 _18105_ (.A1(_08936_),
    .A2(_08937_),
    .A3(_08903_),
    .B1(_08899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08953_));
 sky130_fd_sc_hd__a22oi_2 _18106_ (.A1(_08933_),
    .A2(_08931_),
    .B1(_08900_),
    .B2(_08938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_2 _18107_ (.A(_04259_),
    .B(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08955_));
 sky130_fd_sc_hd__a22oi_2 _18108_ (.A1(\a_l[1] ),
    .A2(\b_l[6] ),
    .B1(\b_l[7] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08956_));
 sky130_fd_sc_hd__a21o_2 _18109_ (.A1(_04259_),
    .A2(_06401_),
    .B1(_08956_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08957_));
 sky130_fd_sc_hd__o21a_2 _18110_ (.A1(_08904_),
    .A2(_08907_),
    .B1(_08909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08958_));
 sky130_fd_sc_hd__o211a_2 _18111_ (.A1(_08904_),
    .A2(_08907_),
    .B1(_08909_),
    .C1(_08957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08959_));
 sky130_fd_sc_hd__nor2_2 _18112_ (.A(_08957_),
    .B(_08958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08960_));
 sky130_fd_sc_hd__nor2_2 _18113_ (.A(_08959_),
    .B(_08960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08961_));
 sky130_fd_sc_hd__or2_2 _18114_ (.A(_08959_),
    .B(_08960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08962_));
 sky130_fd_sc_hd__o2bb2ai_2 _18115_ (.A1_N(_08913_),
    .A2_N(_08929_),
    .B1(_08927_),
    .B2(_08922_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08963_));
 sky130_fd_sc_hd__a21boi_2 _18116_ (.A1(_08913_),
    .A2(_08929_),
    .B1_N(_08928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08964_));
 sky130_fd_sc_hd__nand2_2 _18117_ (.A(\b_l[2] ),
    .B(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_2 _18118_ (.A(\b_l[0] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08966_));
 sky130_fd_sc_hd__nand2_2 _18119_ (.A(\b_l[1] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08967_));
 sky130_fd_sc_hd__a22oi_2 _18120_ (.A1(\b_l[1] ),
    .A2(\a_l[6] ),
    .B1(\a_l[7] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08968_));
 sky130_fd_sc_hd__nand2_2 _18121_ (.A(_08966_),
    .B(_08967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08969_));
 sky130_fd_sc_hd__nand3_2 _18122_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08970_));
 sky130_fd_sc_hd__nand4_2 _18123_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[6] ),
    .D(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08971_));
 sky130_fd_sc_hd__a22oi_2 _18124_ (.A1(\b_l[2] ),
    .A2(\a_l[5] ),
    .B1(_08969_),
    .B2(_08971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08972_));
 sky130_fd_sc_hd__a21bo_2 _18125_ (.A1(_08969_),
    .A2(_08971_),
    .B1_N(_08965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08973_));
 sky130_fd_sc_hd__o2111ai_2 _18126_ (.A1(_09242_),
    .A2(_08970_),
    .B1(\a_l[5] ),
    .C1(_08969_),
    .D1(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08974_));
 sky130_fd_sc_hd__a21o_2 _18127_ (.A1(_08969_),
    .A2(_08971_),
    .B1(_08965_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08975_));
 sky130_fd_sc_hd__o221ai_2 _18128_ (.A1(_09155_),
    .A2(_09210_),
    .B1(_09242_),
    .B2(_08970_),
    .C1(_08969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08976_));
 sky130_fd_sc_hd__nand2_2 _18129_ (.A(_08916_),
    .B(_08921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08977_));
 sky130_fd_sc_hd__o22ai_2 _18130_ (.A1(_04134_),
    .A2(_06681_),
    .B1(_08916_),
    .B2(_08919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08978_));
 sky130_fd_sc_hd__nand2_2 _18131_ (.A(_08920_),
    .B(_08977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08979_));
 sky130_fd_sc_hd__nand3_2 _18132_ (.A(_08975_),
    .B(_08976_),
    .C(_08979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08980_));
 sky130_fd_sc_hd__nand2_2 _18133_ (.A(_08974_),
    .B(_08978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08981_));
 sky130_fd_sc_hd__nand3_2 _18134_ (.A(_08973_),
    .B(_08974_),
    .C(_08978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08982_));
 sky130_fd_sc_hd__nand2_2 _18135_ (.A(\a_l[2] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08983_));
 sky130_fd_sc_hd__nand2_2 _18136_ (.A(\a_l[3] ),
    .B(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08984_));
 sky130_fd_sc_hd__nand2_2 _18137_ (.A(\b_l[3] ),
    .B(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08985_));
 sky130_fd_sc_hd__nand4_2 _18138_ (.A(\a_l[3] ),
    .B(\b_l[3] ),
    .C(\a_l[4] ),
    .D(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08986_));
 sky130_fd_sc_hd__a22oi_2 _18139_ (.A1(\b_l[3] ),
    .A2(\a_l[4] ),
    .B1(\b_l[4] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08987_));
 sky130_fd_sc_hd__nand2_2 _18140_ (.A(_08984_),
    .B(_08985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08988_));
 sky130_fd_sc_hd__a22oi_2 _18141_ (.A1(\a_l[2] ),
    .A2(\b_l[5] ),
    .B1(_08986_),
    .B2(_08988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08989_));
 sky130_fd_sc_hd__and3_2 _18142_ (.A(_08986_),
    .B(\b_l[5] ),
    .C(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08990_));
 sky130_fd_sc_hd__and4_2 _18143_ (.A(_08988_),
    .B(\b_l[5] ),
    .C(\a_l[2] ),
    .D(_08986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08991_));
 sky130_fd_sc_hd__and3_2 _18144_ (.A(_08983_),
    .B(_08986_),
    .C(_08988_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_08992_));
 sky130_fd_sc_hd__a21oi_2 _18145_ (.A1(_08986_),
    .A2(_08988_),
    .B1(_08983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08993_));
 sky130_fd_sc_hd__a21oi_2 _18146_ (.A1(_08990_),
    .A2(_08988_),
    .B1(_08989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08994_));
 sky130_fd_sc_hd__o221ai_2 _18147_ (.A1(_08989_),
    .A2(_08991_),
    .B1(_08972_),
    .B2(_08981_),
    .C1(_08980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08995_));
 sky130_fd_sc_hd__o2bb2ai_2 _18148_ (.A1_N(_08980_),
    .A2_N(_08982_),
    .B1(_08992_),
    .B2(_08993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08996_));
 sky130_fd_sc_hd__o2bb2ai_2 _18149_ (.A1_N(_08980_),
    .A2_N(_08982_),
    .B1(_08989_),
    .B2(_08991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08997_));
 sky130_fd_sc_hd__o211ai_2 _18150_ (.A1(_08992_),
    .A2(_08993_),
    .B1(_08980_),
    .C1(_08982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08998_));
 sky130_fd_sc_hd__a21oi_2 _18151_ (.A1(_08997_),
    .A2(_08998_),
    .B1(_08963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_08999_));
 sky130_fd_sc_hd__nand3_2 _18152_ (.A(_08964_),
    .B(_08995_),
    .C(_08996_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09000_));
 sky130_fd_sc_hd__nand3_2 _18153_ (.A(_08963_),
    .B(_08997_),
    .C(_08998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09001_));
 sky130_fd_sc_hd__nand2_2 _18154_ (.A(_09000_),
    .B(_09001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09002_));
 sky130_fd_sc_hd__and3_2 _18155_ (.A(_09000_),
    .B(_09001_),
    .C(_08961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09003_));
 sky130_fd_sc_hd__nand3_2 _18156_ (.A(_09000_),
    .B(_09001_),
    .C(_08961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09004_));
 sky130_fd_sc_hd__o21ai_2 _18157_ (.A1(_08959_),
    .A2(_08960_),
    .B1(_09002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09005_));
 sky130_fd_sc_hd__a31oi_2 _18158_ (.A1(_08963_),
    .A2(_08997_),
    .A3(_08998_),
    .B1(_08961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09006_));
 sky130_fd_sc_hd__a31o_2 _18159_ (.A1(_08963_),
    .A2(_08997_),
    .A3(_08998_),
    .B1(_08961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09007_));
 sky130_fd_sc_hd__nand2_2 _18160_ (.A(_09006_),
    .B(_09000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09008_));
 sky130_fd_sc_hd__nand2_2 _18161_ (.A(_09002_),
    .B(_08961_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09009_));
 sky130_fd_sc_hd__nand2_2 _18162_ (.A(_08954_),
    .B(_09005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09010_));
 sky130_fd_sc_hd__nand3_2 _18163_ (.A(_09005_),
    .B(_08954_),
    .C(_09004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09011_));
 sky130_fd_sc_hd__o211ai_2 _18164_ (.A1(_08934_),
    .A2(_08953_),
    .B1(_09008_),
    .C1(_09009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09012_));
 sky130_fd_sc_hd__nand2_2 _18165_ (.A(_09011_),
    .B(_09012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09013_));
 sky130_fd_sc_hd__nand3_2 _18166_ (.A(_09011_),
    .B(_09012_),
    .C(_08898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09014_));
 sky130_fd_sc_hd__o2bb2ai_2 _18167_ (.A1_N(_09011_),
    .A2_N(_09012_),
    .B1(_08895_),
    .B2(_08896_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09015_));
 sky130_fd_sc_hd__o221ai_2 _18168_ (.A1(_08895_),
    .A2(_08896_),
    .B1(_09003_),
    .B2(_09010_),
    .C1(_09012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09016_));
 sky130_fd_sc_hd__nand2_2 _18169_ (.A(_09013_),
    .B(_08898_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09017_));
 sky130_fd_sc_hd__nand2_2 _18170_ (.A(_09016_),
    .B(_09017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09018_));
 sky130_fd_sc_hd__and3_2 _18171_ (.A(_09015_),
    .B(_08948_),
    .C(_09014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09019_));
 sky130_fd_sc_hd__nand3_2 _18172_ (.A(_09015_),
    .B(_08948_),
    .C(_09014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09020_));
 sky130_fd_sc_hd__o211ai_2 _18173_ (.A1(_08943_),
    .A2(_08945_),
    .B1(_09016_),
    .C1(_09017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09021_));
 sky130_fd_sc_hd__nand2_2 _18174_ (.A(_09020_),
    .B(_09021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09022_));
 sky130_fd_sc_hd__a2bb2o_2 _18175_ (.A1_N(_08894_),
    .A2_N(_08950_),
    .B1(_09020_),
    .B2(_09021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09023_));
 sky130_fd_sc_hd__o311a_2 _18176_ (.A1(_08894_),
    .A2(_08950_),
    .A3(_09022_),
    .B1(_09023_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00377_));
 sky130_fd_sc_hd__o21ai_2 _18177_ (.A1(_08962_),
    .A2(_08999_),
    .B1(_09001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_2 _18178_ (.A(\a_l[0] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09025_));
 sky130_fd_sc_hd__nand2_2 _18179_ (.A(\a_l[1] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09026_));
 sky130_fd_sc_hd__nand2_2 _18180_ (.A(\a_l[2] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09027_));
 sky130_fd_sc_hd__nand4_2 _18181_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_l[6] ),
    .D(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_2 _18182_ (.A(_09026_),
    .B(_09027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09029_));
 sky130_fd_sc_hd__nand4_2 _18183_ (.A(_09029_),
    .B(\b_l[8] ),
    .C(\a_l[0] ),
    .D(_09028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09030_));
 sky130_fd_sc_hd__nand3_2 _18184_ (.A(_09027_),
    .B(\b_l[7] ),
    .C(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09031_));
 sky130_fd_sc_hd__nand3_2 _18185_ (.A(_09026_),
    .B(\b_l[6] ),
    .C(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09032_));
 sky130_fd_sc_hd__nand3_2 _18186_ (.A(_09025_),
    .B(_09031_),
    .C(_09032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09033_));
 sky130_fd_sc_hd__o21a_2 _18187_ (.A1(_08984_),
    .A2(_08985_),
    .B1(_08983_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09034_));
 sky130_fd_sc_hd__a21oi_2 _18188_ (.A1(_08983_),
    .A2(_08986_),
    .B1(_08987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09035_));
 sky130_fd_sc_hd__a21oi_2 _18189_ (.A1(_09030_),
    .A2(_09033_),
    .B1(_09035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09036_));
 sky130_fd_sc_hd__o2bb2ai_2 _18190_ (.A1_N(_09030_),
    .A2_N(_09033_),
    .B1(_09034_),
    .B2(_08987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09037_));
 sky130_fd_sc_hd__nand3_2 _18191_ (.A(_09030_),
    .B(_09033_),
    .C(_09035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09038_));
 sky130_fd_sc_hd__a22oi_2 _18192_ (.A1(_04259_),
    .A2(_06401_),
    .B1(_09037_),
    .B2(_09038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09039_));
 sky130_fd_sc_hd__a32o_2 _18193_ (.A1(\a_l[1] ),
    .A2(\a_l[0] ),
    .A3(_04259_),
    .B1(_09037_),
    .B2(_09038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09040_));
 sky130_fd_sc_hd__nor2_2 _18194_ (.A(_08955_),
    .B(_09036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09041_));
 sky130_fd_sc_hd__or2_2 _18195_ (.A(_08955_),
    .B(_09036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09042_));
 sky130_fd_sc_hd__nand4_2 _18196_ (.A(_09037_),
    .B(_09038_),
    .C(_04259_),
    .D(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09043_));
 sky130_fd_sc_hd__a21oi_2 _18197_ (.A1(_09041_),
    .A2(_09038_),
    .B1(_09039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09044_));
 sky130_fd_sc_hd__nand2_2 _18198_ (.A(_09040_),
    .B(_09043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09045_));
 sky130_fd_sc_hd__a2bb2oi_2 _18199_ (.A1_N(_08972_),
    .A2_N(_08981_),
    .B1(_08980_),
    .B2(_08994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09046_));
 sky130_fd_sc_hd__o2bb2ai_2 _18200_ (.A1_N(_08994_),
    .A2_N(_08980_),
    .B1(_08972_),
    .B2(_08981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_2 _18201_ (.A(\a_l[3] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09048_));
 sky130_fd_sc_hd__a22oi_2 _18202_ (.A1(\a_l[4] ),
    .A2(\b_l[4] ),
    .B1(\a_l[5] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09049_));
 sky130_fd_sc_hd__nand2_2 _18203_ (.A(\b_l[4] ),
    .B(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09050_));
 sky130_fd_sc_hd__and4_2 _18204_ (.A(\b_l[3] ),
    .B(\a_l[4] ),
    .C(\b_l[4] ),
    .D(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09051_));
 sky130_fd_sc_hd__nand4_2 _18205_ (.A(\b_l[3] ),
    .B(\a_l[4] ),
    .C(\b_l[4] ),
    .D(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09052_));
 sky130_fd_sc_hd__o22a_2 _18206_ (.A1(_09188_),
    .A2(_09220_),
    .B1(_09049_),
    .B2(_09051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09053_));
 sky130_fd_sc_hd__o21ai_2 _18207_ (.A1(_09049_),
    .A2(_09051_),
    .B1(_09048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09054_));
 sky130_fd_sc_hd__a41o_2 _18208_ (.A1(\b_l[3] ),
    .A2(\a_l[4] ),
    .A3(\b_l[4] ),
    .A4(\a_l[5] ),
    .B1(_09048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09055_));
 sky130_fd_sc_hd__nor2_2 _18209_ (.A(_09049_),
    .B(_09055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09056_));
 sky130_fd_sc_hd__o21a_2 _18210_ (.A1(_09049_),
    .A2(_09055_),
    .B1(_09054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09057_));
 sky130_fd_sc_hd__o21ai_2 _18211_ (.A1(_09049_),
    .A2(_09055_),
    .B1(_09054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09058_));
 sky130_fd_sc_hd__nand2_2 _18212_ (.A(_08965_),
    .B(_08971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09059_));
 sky130_fd_sc_hd__o22ai_2 _18213_ (.A1(_09242_),
    .A2(_08970_),
    .B1(_08965_),
    .B2(_08968_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09060_));
 sky130_fd_sc_hd__nand2_2 _18214_ (.A(\b_l[2] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09061_));
 sky130_fd_sc_hd__nand2_2 _18215_ (.A(\b_l[1] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09062_));
 sky130_fd_sc_hd__nand2_2 _18216_ (.A(\b_l[1] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09063_));
 sky130_fd_sc_hd__nand2_2 _18217_ (.A(\b_l[0] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09064_));
 sky130_fd_sc_hd__and4_2 _18218_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[7] ),
    .D(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09065_));
 sky130_fd_sc_hd__nand4_2 _18219_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[7] ),
    .D(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09066_));
 sky130_fd_sc_hd__a22oi_2 _18220_ (.A1(\b_l[1] ),
    .A2(\a_l[7] ),
    .B1(\a_l[8] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09067_));
 sky130_fd_sc_hd__nand2_2 _18221_ (.A(_09063_),
    .B(_09064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09068_));
 sky130_fd_sc_hd__o2bb2ai_2 _18222_ (.A1_N(_09066_),
    .A2_N(_09068_),
    .B1(_09155_),
    .B2(_09231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09069_));
 sky130_fd_sc_hd__o2111ai_2 _18223_ (.A1(_04134_),
    .A2(_06867_),
    .B1(\b_l[2] ),
    .C1(\a_l[6] ),
    .D1(_09068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09070_));
 sky130_fd_sc_hd__a21oi_2 _18224_ (.A1(_09066_),
    .A2(_09068_),
    .B1(_09061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_2 _18225_ (.A(_09061_),
    .B(_09066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09072_));
 sky130_fd_sc_hd__o2bb2ai_2 _18226_ (.A1_N(_08969_),
    .A2_N(_09059_),
    .B1(_09067_),
    .B2(_09072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09073_));
 sky130_fd_sc_hd__nand3_2 _18227_ (.A(_09069_),
    .B(_09070_),
    .C(_09060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09074_));
 sky130_fd_sc_hd__o21ai_2 _18228_ (.A1(_09071_),
    .A2(_09073_),
    .B1(_09074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09075_));
 sky130_fd_sc_hd__o221ai_2 _18229_ (.A1(_09071_),
    .A2(_09073_),
    .B1(_09053_),
    .B2(_09056_),
    .C1(_09074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09076_));
 sky130_fd_sc_hd__nand2_2 _18230_ (.A(_09075_),
    .B(_09057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09077_));
 sky130_fd_sc_hd__o211ai_2 _18231_ (.A1(_09071_),
    .A2(_09073_),
    .B1(_09074_),
    .C1(_09057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09078_));
 sky130_fd_sc_hd__o21ai_2 _18232_ (.A1(_09053_),
    .A2(_09056_),
    .B1(_09075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09079_));
 sky130_fd_sc_hd__a31o_2 _18233_ (.A1(_08973_),
    .A2(_08974_),
    .A3(_08978_),
    .B1(_08994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09080_));
 sky130_fd_sc_hd__a21boi_2 _18234_ (.A1(_09058_),
    .A2(_09075_),
    .B1_N(_08980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09081_));
 sky130_fd_sc_hd__nand3_2 _18235_ (.A(_09047_),
    .B(_09078_),
    .C(_09079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09082_));
 sky130_fd_sc_hd__nand3_2 _18236_ (.A(_09077_),
    .B(_09046_),
    .C(_09076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09083_));
 sky130_fd_sc_hd__nand2_2 _18237_ (.A(_09082_),
    .B(_09083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09084_));
 sky130_fd_sc_hd__nand3_2 _18238_ (.A(_09045_),
    .B(_09082_),
    .C(_09083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09085_));
 sky130_fd_sc_hd__nand2_2 _18239_ (.A(_09084_),
    .B(_09044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09086_));
 sky130_fd_sc_hd__o211ai_2 _18240_ (.A1(_08999_),
    .A2(_09006_),
    .B1(_09085_),
    .C1(_09086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09087_));
 sky130_fd_sc_hd__nand3_2 _18241_ (.A(_09082_),
    .B(_09083_),
    .C(_09044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09088_));
 sky130_fd_sc_hd__a21oi_2 _18242_ (.A1(_09082_),
    .A2(_09083_),
    .B1(_09044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09089_));
 sky130_fd_sc_hd__a22o_2 _18243_ (.A1(_09040_),
    .A2(_09043_),
    .B1(_09082_),
    .B2(_09083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09090_));
 sky130_fd_sc_hd__nand3_2 _18244_ (.A(_09000_),
    .B(_09007_),
    .C(_09088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09091_));
 sky130_fd_sc_hd__nand3_2 _18245_ (.A(_09090_),
    .B(_09024_),
    .C(_09088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09092_));
 sky130_fd_sc_hd__o2bb2ai_2 _18246_ (.A1_N(_09087_),
    .A2_N(_09092_),
    .B1(_08957_),
    .B2(_08958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09093_));
 sky130_fd_sc_hd__o211ai_2 _18247_ (.A1(_09089_),
    .A2(_09091_),
    .B1(_08960_),
    .C1(_09087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09094_));
 sky130_fd_sc_hd__o2bb2ai_2 _18248_ (.A1_N(_08898_),
    .A2_N(_09012_),
    .B1(_09003_),
    .B2(_09010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09095_));
 sky130_fd_sc_hd__a21oi_2 _18249_ (.A1(_09093_),
    .A2(_09094_),
    .B1(_09095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09096_));
 sky130_fd_sc_hd__a21o_2 _18250_ (.A1(_09093_),
    .A2(_09094_),
    .B1(_09095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09097_));
 sky130_fd_sc_hd__nand2_2 _18251_ (.A(_09019_),
    .B(_09097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09098_));
 sky130_fd_sc_hd__nand3_2 _18252_ (.A(_09093_),
    .B(_09095_),
    .C(_09094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09099_));
 sky130_fd_sc_hd__nand2_2 _18253_ (.A(_09097_),
    .B(_09099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09100_));
 sky130_fd_sc_hd__a21boi_2 _18254_ (.A1(_09021_),
    .A2(_08951_),
    .B1_N(_09020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09101_));
 sky130_fd_sc_hd__and2_2 _18255_ (.A(_09101_),
    .B(_09100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09102_));
 sky130_fd_sc_hd__and4_2 _18256_ (.A(_09097_),
    .B(_08951_),
    .C(_09021_),
    .D(_09099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09103_));
 sky130_fd_sc_hd__o2111ai_2 _18257_ (.A1(_08948_),
    .A2(_09018_),
    .B1(_08951_),
    .C1(_09099_),
    .D1(_09097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09104_));
 sky130_fd_sc_hd__a31o_2 _18258_ (.A1(_08948_),
    .A2(_09018_),
    .A3(_09097_),
    .B1(_09103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09105_));
 sky130_fd_sc_hd__or4b_2 _18259_ (.A(_08856_),
    .B(_08890_),
    .C(_08950_),
    .D_N(_09018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09106_));
 sky130_fd_sc_hd__nand4_2 _18260_ (.A(_08892_),
    .B(_08947_),
    .C(_08949_),
    .D(_09018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09107_));
 sky130_fd_sc_hd__o21a_2 _18261_ (.A1(_09105_),
    .A2(_09102_),
    .B1(_09106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09108_));
 sky130_fd_sc_hd__a21oi_2 _18262_ (.A1(_09101_),
    .A2(_09100_),
    .B1(_09107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09109_));
 sky130_fd_sc_hd__nor3_2 _18263_ (.A(rst),
    .B(_09108_),
    .C(_09109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00378_));
 sky130_fd_sc_hd__a31o_2 _18264_ (.A1(_09090_),
    .A2(_09024_),
    .A3(_09088_),
    .B1(_08960_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09110_));
 sky130_fd_sc_hd__o2bb2ai_2 _18265_ (.A1_N(_08960_),
    .A2_N(_09087_),
    .B1(_09089_),
    .B2(_09091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09111_));
 sky130_fd_sc_hd__a2bb2oi_2 _18266_ (.A1_N(_09089_),
    .A2_N(_09091_),
    .B1(_08960_),
    .B2(_09087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09112_));
 sky130_fd_sc_hd__o21ai_2 _18267_ (.A1(_04260_),
    .A2(_06441_),
    .B1(_09030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09113_));
 sky130_fd_sc_hd__a21oi_2 _18268_ (.A1(_09048_),
    .A2(_09052_),
    .B1(_09049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09114_));
 sky130_fd_sc_hd__nand2_2 _18269_ (.A(\a_l[1] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09115_));
 sky130_fd_sc_hd__nand2_2 _18270_ (.A(\a_l[2] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09116_));
 sky130_fd_sc_hd__nand2_2 _18271_ (.A(\a_l[3] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09117_));
 sky130_fd_sc_hd__nand4_2 _18272_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_l[6] ),
    .D(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09118_));
 sky130_fd_sc_hd__nand2_2 _18273_ (.A(_09116_),
    .B(_09117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09119_));
 sky130_fd_sc_hd__nand3_2 _18274_ (.A(_09116_),
    .B(\b_l[6] ),
    .C(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09120_));
 sky130_fd_sc_hd__nand3_2 _18275_ (.A(_09117_),
    .B(\b_l[7] ),
    .C(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09121_));
 sky130_fd_sc_hd__nand3_2 _18276_ (.A(_09115_),
    .B(_09120_),
    .C(_09121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09122_));
 sky130_fd_sc_hd__nand4_2 _18277_ (.A(_09119_),
    .B(\b_l[8] ),
    .C(\a_l[1] ),
    .D(_09118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09123_));
 sky130_fd_sc_hd__nand3_2 _18278_ (.A(_09114_),
    .B(_09122_),
    .C(_09123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09124_));
 sky130_fd_sc_hd__a21o_2 _18279_ (.A1(_09122_),
    .A2(_09123_),
    .B1(_09114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09125_));
 sky130_fd_sc_hd__a21oi_2 _18280_ (.A1(_09124_),
    .A2(_09125_),
    .B1(_09113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09126_));
 sky130_fd_sc_hd__and3_2 _18281_ (.A(_09113_),
    .B(_09124_),
    .C(_09125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09127_));
 sky130_fd_sc_hd__nand3_2 _18282_ (.A(_09113_),
    .B(_09124_),
    .C(_09125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09128_));
 sky130_fd_sc_hd__o2111ai_2 _18283_ (.A1(_04260_),
    .A2(_06441_),
    .B1(_09030_),
    .C1(_09124_),
    .D1(_09125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09129_));
 sky130_fd_sc_hd__a22o_2 _18284_ (.A1(_09028_),
    .A2(_09030_),
    .B1(_09124_),
    .B2(_09125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09130_));
 sky130_fd_sc_hd__nand2_2 _18285_ (.A(_09129_),
    .B(_09130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09131_));
 sky130_fd_sc_hd__o2bb2ai_2 _18286_ (.A1_N(_09058_),
    .A2_N(_09074_),
    .B1(_09073_),
    .B2(_09071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09132_));
 sky130_fd_sc_hd__a2bb2oi_2 _18287_ (.A1_N(_09071_),
    .A2_N(_09073_),
    .B1(_09074_),
    .B2(_09058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09133_));
 sky130_fd_sc_hd__nand2_2 _18288_ (.A(\a_l[4] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09134_));
 sky130_fd_sc_hd__nand2_2 _18289_ (.A(\b_l[3] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09135_));
 sky130_fd_sc_hd__nand4_2 _18290_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[5] ),
    .D(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09136_));
 sky130_fd_sc_hd__a22oi_2 _18291_ (.A1(\b_l[4] ),
    .A2(\a_l[5] ),
    .B1(\a_l[6] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09137_));
 sky130_fd_sc_hd__nand2_2 _18292_ (.A(_09050_),
    .B(_09135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09138_));
 sky130_fd_sc_hd__o21a_2 _18293_ (.A1(_04182_),
    .A2(_06681_),
    .B1(_09134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09139_));
 sky130_fd_sc_hd__o221a_2 _18294_ (.A1(_09199_),
    .A2(_09220_),
    .B1(_04182_),
    .B2(_06681_),
    .C1(_09138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09140_));
 sky130_fd_sc_hd__a21oi_2 _18295_ (.A1(_09136_),
    .A2(_09138_),
    .B1(_09134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09141_));
 sky130_fd_sc_hd__o2bb2ai_2 _18296_ (.A1_N(_09136_),
    .A2_N(_09138_),
    .B1(_09199_),
    .B2(_09220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09142_));
 sky130_fd_sc_hd__a41o_2 _18297_ (.A1(\b_l[3] ),
    .A2(\b_l[4] ),
    .A3(\a_l[5] ),
    .A4(\a_l[6] ),
    .B1(_09134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09143_));
 sky130_fd_sc_hd__o21ai_2 _18298_ (.A1(_09137_),
    .A2(_09143_),
    .B1(_09142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09145_));
 sky130_fd_sc_hd__a21oi_2 _18299_ (.A1(_09063_),
    .A2(_09064_),
    .B1(_09061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09146_));
 sky130_fd_sc_hd__nand2_2 _18300_ (.A(_09068_),
    .B(_09072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09147_));
 sky130_fd_sc_hd__nand2_2 _18301_ (.A(\b_l[0] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09148_));
 sky130_fd_sc_hd__a22oi_2 _18302_ (.A1(\b_l[1] ),
    .A2(\a_l[8] ),
    .B1(\a_l[9] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09149_));
 sky130_fd_sc_hd__nand2_2 _18303_ (.A(_09062_),
    .B(_09148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09150_));
 sky130_fd_sc_hd__nand4_2 _18304_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[8] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_2 _18305_ (.A(_09150_),
    .B(_09151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09152_));
 sky130_fd_sc_hd__nor2_2 _18306_ (.A(_09155_),
    .B(_09242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_2 _18307_ (.A(\b_l[2] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09154_));
 sky130_fd_sc_hd__nand2_2 _18308_ (.A(_09152_),
    .B(_09153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09156_));
 sky130_fd_sc_hd__o211ai_2 _18309_ (.A1(_09155_),
    .A2(_09242_),
    .B1(_09150_),
    .C1(_09151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09157_));
 sky130_fd_sc_hd__nand4_2 _18310_ (.A(_09150_),
    .B(_09151_),
    .C(\b_l[2] ),
    .D(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09158_));
 sky130_fd_sc_hd__o2bb2ai_2 _18311_ (.A1_N(_09150_),
    .A2_N(_09151_),
    .B1(_09155_),
    .B2(_09242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09159_));
 sky130_fd_sc_hd__o211a_2 _18312_ (.A1(_09065_),
    .A2(_09146_),
    .B1(_09158_),
    .C1(_09159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09160_));
 sky130_fd_sc_hd__o211ai_2 _18313_ (.A1(_09065_),
    .A2(_09146_),
    .B1(_09158_),
    .C1(_09159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09161_));
 sky130_fd_sc_hd__nand3_2 _18314_ (.A(_09156_),
    .B(_09157_),
    .C(_09147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09162_));
 sky130_fd_sc_hd__nand2_2 _18315_ (.A(_09161_),
    .B(_09162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09163_));
 sky130_fd_sc_hd__o21ai_2 _18316_ (.A1(_09140_),
    .A2(_09141_),
    .B1(_09162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09164_));
 sky130_fd_sc_hd__nand2_2 _18317_ (.A(_09163_),
    .B(_09145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09165_));
 sky130_fd_sc_hd__nand3_2 _18318_ (.A(_09161_),
    .B(_09162_),
    .C(_09145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09167_));
 sky130_fd_sc_hd__o21ai_2 _18319_ (.A1(_09140_),
    .A2(_09141_),
    .B1(_09163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09168_));
 sky130_fd_sc_hd__o211a_2 _18320_ (.A1(_09164_),
    .A2(_09160_),
    .B1(_09133_),
    .C1(_09165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09169_));
 sky130_fd_sc_hd__o211ai_2 _18321_ (.A1(_09164_),
    .A2(_09160_),
    .B1(_09133_),
    .C1(_09165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09170_));
 sky130_fd_sc_hd__nand3_2 _18322_ (.A(_09168_),
    .B(_09132_),
    .C(_09167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_2 _18323_ (.A(_09170_),
    .B(_09171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09172_));
 sky130_fd_sc_hd__o21ai_2 _18324_ (.A1(_09126_),
    .A2(_09127_),
    .B1(_09172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09173_));
 sky130_fd_sc_hd__nand3_2 _18325_ (.A(_09131_),
    .B(_09170_),
    .C(_09171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09174_));
 sky130_fd_sc_hd__o21ai_2 _18326_ (.A1(_09126_),
    .A2(_09127_),
    .B1(_09171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09175_));
 sky130_fd_sc_hd__o211ai_2 _18327_ (.A1(_09126_),
    .A2(_09127_),
    .B1(_09170_),
    .C1(_09171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09176_));
 sky130_fd_sc_hd__nand2_2 _18328_ (.A(_09172_),
    .B(_09131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09178_));
 sky130_fd_sc_hd__nand2_2 _18329_ (.A(_09045_),
    .B(_09082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09179_));
 sky130_fd_sc_hd__a32oi_2 _18330_ (.A1(_09081_),
    .A2(_09080_),
    .A3(_09078_),
    .B1(_09083_),
    .B2(_09044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09180_));
 sky130_fd_sc_hd__a21boi_2 _18331_ (.A1(_09045_),
    .A2(_09082_),
    .B1_N(_09083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09181_));
 sky130_fd_sc_hd__nand3_2 _18332_ (.A(_09173_),
    .B(_09174_),
    .C(_09181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09182_));
 sky130_fd_sc_hd__a22oi_2 _18333_ (.A1(_09172_),
    .A2(_09131_),
    .B1(_09083_),
    .B2(_09179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09183_));
 sky130_fd_sc_hd__and3_2 _18334_ (.A(_09176_),
    .B(_09178_),
    .C(_09180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09184_));
 sky130_fd_sc_hd__o211ai_2 _18335_ (.A1(_09169_),
    .A2(_09175_),
    .B1(_09180_),
    .C1(_09178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09185_));
 sky130_fd_sc_hd__nand2_2 _18336_ (.A(_09182_),
    .B(_09185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09186_));
 sky130_fd_sc_hd__nand2_2 _18337_ (.A(\a_l[0] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09187_));
 sky130_fd_sc_hd__o31a_2 _18338_ (.A1(_04260_),
    .A2(_06402_),
    .A3(_09036_),
    .B1(_09038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09189_));
 sky130_fd_sc_hd__a21oi_2 _18339_ (.A1(_09038_),
    .A2(_09042_),
    .B1(_09187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09190_));
 sky130_fd_sc_hd__a21o_2 _18340_ (.A1(_09038_),
    .A2(_09042_),
    .B1(_09187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09191_));
 sky130_fd_sc_hd__o311a_2 _18341_ (.A1(_04260_),
    .A2(_06402_),
    .A3(_09036_),
    .B1(_09038_),
    .C1(_09187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09192_));
 sky130_fd_sc_hd__nand2_2 _18342_ (.A(_09187_),
    .B(_09189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09193_));
 sky130_fd_sc_hd__nor2_2 _18343_ (.A(_09190_),
    .B(_09192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_2 _18344_ (.A(_09191_),
    .B(_09193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09195_));
 sky130_fd_sc_hd__nand2_2 _18345_ (.A(_09186_),
    .B(_09194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09196_));
 sky130_fd_sc_hd__o211ai_2 _18346_ (.A1(_09190_),
    .A2(_09192_),
    .B1(_09182_),
    .C1(_09185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09197_));
 sky130_fd_sc_hd__o2bb2ai_2 _18347_ (.A1_N(_09182_),
    .A2_N(_09185_),
    .B1(_09190_),
    .B2(_09192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09198_));
 sky130_fd_sc_hd__nand4_2 _18348_ (.A(_09182_),
    .B(_09185_),
    .C(_09191_),
    .D(_09193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09200_));
 sky130_fd_sc_hd__a22oi_2 _18349_ (.A1(_09087_),
    .A2(_09110_),
    .B1(_09198_),
    .B2(_09200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09201_));
 sky130_fd_sc_hd__nand3_2 _18350_ (.A(_09112_),
    .B(_09196_),
    .C(_09197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09202_));
 sky130_fd_sc_hd__a21oi_2 _18351_ (.A1(_09186_),
    .A2(_09195_),
    .B1(_09112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09203_));
 sky130_fd_sc_hd__nand3_2 _18352_ (.A(_09198_),
    .B(_09200_),
    .C(_09111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09204_));
 sky130_fd_sc_hd__inv_2 _18353_ (.A(_09204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09205_));
 sky130_fd_sc_hd__a21boi_2 _18354_ (.A1(_09202_),
    .A2(_09204_),
    .B1_N(_09099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09206_));
 sky130_fd_sc_hd__a211oi_2 _18355_ (.A1(_09203_),
    .A2(_09200_),
    .B1(_09099_),
    .C1(_09201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09207_));
 sky130_fd_sc_hd__o22ai_2 _18356_ (.A1(_09020_),
    .A2(_09096_),
    .B1(_09206_),
    .B2(_09207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09208_));
 sky130_fd_sc_hd__o31a_2 _18357_ (.A1(_09020_),
    .A2(_09096_),
    .A3(_09206_),
    .B1(_09208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09209_));
 sky130_fd_sc_hd__o21ai_2 _18358_ (.A1(_09106_),
    .A2(_09102_),
    .B1(_09104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09211_));
 sky130_fd_sc_hd__o31a_2 _18359_ (.A1(_09103_),
    .A2(_09109_),
    .A3(_09209_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09212_));
 sky130_fd_sc_hd__a21boi_2 _18360_ (.A1(_09209_),
    .A2(_09211_),
    .B1_N(_09212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00379_));
 sky130_fd_sc_hd__a31oi_2 _18361_ (.A1(_09173_),
    .A2(_09174_),
    .A3(_09181_),
    .B1(_09194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09213_));
 sky130_fd_sc_hd__a31o_2 _18362_ (.A1(_09173_),
    .A2(_09174_),
    .A3(_09181_),
    .B1(_09194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09214_));
 sky130_fd_sc_hd__a22oi_2 _18363_ (.A1(_09183_),
    .A2(_09176_),
    .B1(_09182_),
    .B2(_09195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09215_));
 sky130_fd_sc_hd__nand2_2 _18364_ (.A(\a_l[1] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09216_));
 sky130_fd_sc_hd__and3_2 _18365_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .C(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09217_));
 sky130_fd_sc_hd__a22oi_2 _18366_ (.A1(\a_l[1] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09218_));
 sky130_fd_sc_hd__a31o_2 _18367_ (.A1(\b_l[9] ),
    .A2(\b_l[10] ),
    .A3(_06401_),
    .B1(_09218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09219_));
 sky130_fd_sc_hd__a31o_2 _18368_ (.A1(_09114_),
    .A2(_09122_),
    .A3(_09123_),
    .B1(_09127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09221_));
 sky130_fd_sc_hd__inv_2 _18369_ (.A(_09221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09222_));
 sky130_fd_sc_hd__a21oi_2 _18370_ (.A1(_09124_),
    .A2(_09128_),
    .B1(_09219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09223_));
 sky130_fd_sc_hd__and3_2 _18371_ (.A(_09124_),
    .B(_09128_),
    .C(_09219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09224_));
 sky130_fd_sc_hd__nor2_2 _18372_ (.A(_09223_),
    .B(_09224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09225_));
 sky130_fd_sc_hd__o21ai_2 _18373_ (.A1(_09126_),
    .A2(_09127_),
    .B1(_09170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09226_));
 sky130_fd_sc_hd__a21oi_2 _18374_ (.A1(_09131_),
    .A2(_09171_),
    .B1(_09169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09227_));
 sky130_fd_sc_hd__nand2_2 _18375_ (.A(_09161_),
    .B(_09145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09228_));
 sky130_fd_sc_hd__nand2_2 _18376_ (.A(_09161_),
    .B(_09164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09229_));
 sky130_fd_sc_hd__nand2_2 _18377_ (.A(_09162_),
    .B(_09228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09230_));
 sky130_fd_sc_hd__a21o_2 _18378_ (.A1(_09151_),
    .A2(_09154_),
    .B1(_09149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09232_));
 sky130_fd_sc_hd__a21oi_2 _18379_ (.A1(_09151_),
    .A2(_09154_),
    .B1(_09149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2_2 _18380_ (.A(\b_l[2] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09234_));
 sky130_fd_sc_hd__nand2_2 _18381_ (.A(\b_l[1] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_2 _18382_ (.A(\b_l[0] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09236_));
 sky130_fd_sc_hd__a22oi_2 _18383_ (.A1(\b_l[1] ),
    .A2(\a_l[9] ),
    .B1(\a_l[10] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09237_));
 sky130_fd_sc_hd__nand2_2 _18384_ (.A(_09235_),
    .B(_09236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09238_));
 sky130_fd_sc_hd__nand4_2 _18385_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[9] ),
    .D(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09239_));
 sky130_fd_sc_hd__o2bb2ai_2 _18386_ (.A1_N(_09238_),
    .A2_N(_09239_),
    .B1(_09155_),
    .B2(_09253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09240_));
 sky130_fd_sc_hd__o2111ai_2 _18387_ (.A1(_04134_),
    .A2(_07100_),
    .B1(\b_l[2] ),
    .C1(\a_l[8] ),
    .D1(_09238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09241_));
 sky130_fd_sc_hd__nand3_2 _18388_ (.A(_09233_),
    .B(_09240_),
    .C(_09241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09243_));
 sky130_fd_sc_hd__a21o_2 _18389_ (.A1(_09238_),
    .A2(_09239_),
    .B1(_09234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09244_));
 sky130_fd_sc_hd__o221ai_2 _18390_ (.A1(_09155_),
    .A2(_09253_),
    .B1(_04134_),
    .B2(_07100_),
    .C1(_09238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09245_));
 sky130_fd_sc_hd__and3_2 _18391_ (.A(_09244_),
    .B(_09245_),
    .C(_09232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09246_));
 sky130_fd_sc_hd__nand3_2 _18392_ (.A(_09244_),
    .B(_09245_),
    .C(_09232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09247_));
 sky130_fd_sc_hd__nand2_2 _18393_ (.A(\a_l[5] ),
    .B(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09248_));
 sky130_fd_sc_hd__a22oi_2 _18394_ (.A1(\b_l[4] ),
    .A2(\a_l[6] ),
    .B1(\a_l[7] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09249_));
 sky130_fd_sc_hd__a22o_2 _18395_ (.A1(\b_l[4] ),
    .A2(\a_l[6] ),
    .B1(\a_l[7] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09250_));
 sky130_fd_sc_hd__nand4_2 _18396_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[6] ),
    .D(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09251_));
 sky130_fd_sc_hd__o2bb2a_2 _18397_ (.A1_N(_09250_),
    .A2_N(_09251_),
    .B1(_09210_),
    .B2(_09220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09252_));
 sky130_fd_sc_hd__a22o_2 _18398_ (.A1(\a_l[5] ),
    .A2(\b_l[5] ),
    .B1(_09250_),
    .B2(_09251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09254_));
 sky130_fd_sc_hd__and4_2 _18399_ (.A(_09250_),
    .B(_09251_),
    .C(\a_l[5] ),
    .D(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09255_));
 sky130_fd_sc_hd__nand4_2 _18400_ (.A(_09250_),
    .B(_09251_),
    .C(\a_l[5] ),
    .D(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09256_));
 sky130_fd_sc_hd__a21oi_2 _18401_ (.A1(_09250_),
    .A2(_09251_),
    .B1(_09248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09257_));
 sky130_fd_sc_hd__o311a_2 _18402_ (.A1(_09231_),
    .A2(_09242_),
    .A3(_04182_),
    .B1(_09248_),
    .C1(_09250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09258_));
 sky130_fd_sc_hd__nand2_2 _18403_ (.A(_09254_),
    .B(_09256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09259_));
 sky130_fd_sc_hd__nand3_2 _18404_ (.A(_09243_),
    .B(_09247_),
    .C(_09259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09260_));
 sky130_fd_sc_hd__o2bb2ai_2 _18405_ (.A1_N(_09243_),
    .A2_N(_09247_),
    .B1(_09257_),
    .B2(_09258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09261_));
 sky130_fd_sc_hd__o2bb2ai_2 _18406_ (.A1_N(_09243_),
    .A2_N(_09247_),
    .B1(_09252_),
    .B2(_09255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09262_));
 sky130_fd_sc_hd__o211ai_2 _18407_ (.A1(_09257_),
    .A2(_09258_),
    .B1(_09243_),
    .C1(_09247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09263_));
 sky130_fd_sc_hd__nand3_2 _18408_ (.A(_09230_),
    .B(_09260_),
    .C(_09261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09265_));
 sky130_fd_sc_hd__nand3_2 _18409_ (.A(_09229_),
    .B(_09262_),
    .C(_09263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09266_));
 sky130_fd_sc_hd__o31a_2 _18410_ (.A1(_09144_),
    .A2(_09188_),
    .A3(_04260_),
    .B1(_09123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09267_));
 sky130_fd_sc_hd__o21ai_2 _18411_ (.A1(_09134_),
    .A2(_09137_),
    .B1(_09136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09268_));
 sky130_fd_sc_hd__and2_2 _18412_ (.A(\a_l[2] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09269_));
 sky130_fd_sc_hd__nand2_2 _18413_ (.A(\a_l[2] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09270_));
 sky130_fd_sc_hd__nand2_2 _18414_ (.A(\a_l[3] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09271_));
 sky130_fd_sc_hd__nand2_2 _18415_ (.A(\a_l[4] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09272_));
 sky130_fd_sc_hd__a22oi_2 _18416_ (.A1(\a_l[4] ),
    .A2(\b_l[6] ),
    .B1(\b_l[7] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09273_));
 sky130_fd_sc_hd__nand2_2 _18417_ (.A(_09271_),
    .B(_09272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09274_));
 sky130_fd_sc_hd__nand4_2 _18418_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_l[6] ),
    .D(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09276_));
 sky130_fd_sc_hd__o221ai_2 _18419_ (.A1(_09144_),
    .A2(_09264_),
    .B1(_04260_),
    .B2(_06521_),
    .C1(_09274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09277_));
 sky130_fd_sc_hd__a21o_2 _18420_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09278_));
 sky130_fd_sc_hd__a21o_2 _18421_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09279_));
 sky130_fd_sc_hd__o2111ai_2 _18422_ (.A1(_04260_),
    .A2(_06521_),
    .B1(\a_l[2] ),
    .C1(\b_l[8] ),
    .D1(_09274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09280_));
 sky130_fd_sc_hd__o211a_2 _18423_ (.A1(_09137_),
    .A2(_09139_),
    .B1(_09277_),
    .C1(_09278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09281_));
 sky130_fd_sc_hd__o211ai_2 _18424_ (.A1(_09137_),
    .A2(_09139_),
    .B1(_09277_),
    .C1(_09278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3_2 _18425_ (.A(_09279_),
    .B(_09280_),
    .C(_09268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09283_));
 sky130_fd_sc_hd__a21oi_2 _18426_ (.A1(_09282_),
    .A2(_09283_),
    .B1(_09267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09284_));
 sky130_fd_sc_hd__a21o_2 _18427_ (.A1(_09282_),
    .A2(_09283_),
    .B1(_09267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09285_));
 sky130_fd_sc_hd__and3_2 _18428_ (.A(_09282_),
    .B(_09283_),
    .C(_09267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09287_));
 sky130_fd_sc_hd__o2111ai_2 _18429_ (.A1(_04260_),
    .A2(_06480_),
    .B1(_09123_),
    .C1(_09282_),
    .D1(_09283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09288_));
 sky130_fd_sc_hd__nand2_2 _18430_ (.A(_09285_),
    .B(_09288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09289_));
 sky130_fd_sc_hd__a21oi_2 _18431_ (.A1(_09265_),
    .A2(_09266_),
    .B1(_09289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_2 _18432_ (.A(_09265_),
    .B(_09289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09291_));
 sky130_fd_sc_hd__nand3_2 _18433_ (.A(_09265_),
    .B(_09266_),
    .C(_09289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09292_));
 sky130_fd_sc_hd__nand4_2 _18434_ (.A(_09265_),
    .B(_09266_),
    .C(_09285_),
    .D(_09288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09293_));
 sky130_fd_sc_hd__o2bb2ai_2 _18435_ (.A1_N(_09265_),
    .A2_N(_09266_),
    .B1(_09284_),
    .B2(_09287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09294_));
 sky130_fd_sc_hd__nand3_2 _18436_ (.A(_09171_),
    .B(_09226_),
    .C(_09292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09295_));
 sky130_fd_sc_hd__nand3_2 _18437_ (.A(_09227_),
    .B(_09293_),
    .C(_09294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09296_));
 sky130_fd_sc_hd__o21ai_2 _18438_ (.A1(_09290_),
    .A2(_09295_),
    .B1(_09296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09298_));
 sky130_fd_sc_hd__o221ai_2 _18439_ (.A1(_09223_),
    .A2(_09224_),
    .B1(_09290_),
    .B2(_09295_),
    .C1(_09296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_2 _18440_ (.A(_09298_),
    .B(_09225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09300_));
 sky130_fd_sc_hd__o211ai_2 _18441_ (.A1(_09290_),
    .A2(_09295_),
    .B1(_09225_),
    .C1(_09296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09301_));
 sky130_fd_sc_hd__o21ai_2 _18442_ (.A1(_09223_),
    .A2(_09224_),
    .B1(_09298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09302_));
 sky130_fd_sc_hd__a22oi_2 _18443_ (.A1(_09298_),
    .A2(_09225_),
    .B1(_09214_),
    .B2(_09185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09303_));
 sky130_fd_sc_hd__o211ai_2 _18444_ (.A1(_09184_),
    .A2(_09213_),
    .B1(_09299_),
    .C1(_09300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09304_));
 sky130_fd_sc_hd__and3_2 _18445_ (.A(_09302_),
    .B(_09215_),
    .C(_09301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09305_));
 sky130_fd_sc_hd__nand3_2 _18446_ (.A(_09302_),
    .B(_09215_),
    .C(_09301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09306_));
 sky130_fd_sc_hd__o2bb2ai_2 _18447_ (.A1_N(_09304_),
    .A2_N(_09306_),
    .B1(_09187_),
    .B2(_09189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_2 _18448_ (.A(_09304_),
    .B(_09190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09309_));
 sky130_fd_sc_hd__o211ai_2 _18449_ (.A1(_09187_),
    .A2(_09189_),
    .B1(_09304_),
    .C1(_09306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09310_));
 sky130_fd_sc_hd__a21o_2 _18450_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_09191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09311_));
 sky130_fd_sc_hd__nand3_2 _18451_ (.A(_09204_),
    .B(_09310_),
    .C(_09311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09312_));
 sky130_fd_sc_hd__o211a_2 _18452_ (.A1(_09305_),
    .A2(_09309_),
    .B1(_09205_),
    .C1(_09307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09313_));
 sky130_fd_sc_hd__o211ai_2 _18453_ (.A1(_09305_),
    .A2(_09309_),
    .B1(_09205_),
    .C1(_09307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09314_));
 sky130_fd_sc_hd__a21oi_2 _18454_ (.A1(_09312_),
    .A2(_09314_),
    .B1(_09207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09315_));
 sky130_fd_sc_hd__a21o_2 _18455_ (.A1(_09207_),
    .A2(_09312_),
    .B1(_09315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09316_));
 sky130_fd_sc_hd__a21oi_2 _18456_ (.A1(_09202_),
    .A2(_09204_),
    .B1(_09019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09317_));
 sky130_fd_sc_hd__o22ai_2 _18457_ (.A1(_09098_),
    .A2(_09206_),
    .B1(_09317_),
    .B2(_09104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09318_));
 sky130_fd_sc_hd__a21oi_2 _18458_ (.A1(_09208_),
    .A2(_09109_),
    .B1(_09318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09320_));
 sky130_fd_sc_hd__a21oi_2 _18459_ (.A1(_09316_),
    .A2(_09320_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09321_));
 sky130_fd_sc_hd__o21a_2 _18460_ (.A1(_09315_),
    .A2(_09320_),
    .B1(_09321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00380_));
 sky130_fd_sc_hd__o2bb2a_2 _18461_ (.A1_N(_09207_),
    .A2_N(_09312_),
    .B1(_09315_),
    .B2(_09320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09322_));
 sky130_fd_sc_hd__o2bb2ai_2 _18462_ (.A1_N(_09225_),
    .A2_N(_09296_),
    .B1(_09295_),
    .B2(_09290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09323_));
 sky130_fd_sc_hd__a2bb2oi_2 _18463_ (.A1_N(_09290_),
    .A2_N(_09295_),
    .B1(_09225_),
    .B2(_09296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09324_));
 sky130_fd_sc_hd__nand2_2 _18464_ (.A(_09266_),
    .B(_09291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09325_));
 sky130_fd_sc_hd__a21boi_2 _18465_ (.A1(_09265_),
    .A2(_09289_),
    .B1_N(_09266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09326_));
 sky130_fd_sc_hd__o21ai_2 _18466_ (.A1(_09248_),
    .A2(_09249_),
    .B1(_09251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09327_));
 sky130_fd_sc_hd__o21a_2 _18467_ (.A1(_09248_),
    .A2(_09249_),
    .B1(_09251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09328_));
 sky130_fd_sc_hd__nand2_2 _18468_ (.A(\a_l[3] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09330_));
 sky130_fd_sc_hd__nand2_2 _18469_ (.A(\a_l[4] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09331_));
 sky130_fd_sc_hd__nand2_2 _18470_ (.A(\a_l[5] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09332_));
 sky130_fd_sc_hd__a22oi_2 _18471_ (.A1(\a_l[5] ),
    .A2(\b_l[6] ),
    .B1(\b_l[7] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_2 _18472_ (.A(_09331_),
    .B(_09332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09334_));
 sky130_fd_sc_hd__nand4_2 _18473_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_l[6] ),
    .D(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09335_));
 sky130_fd_sc_hd__a41o_2 _18474_ (.A1(\a_l[4] ),
    .A2(\a_l[5] ),
    .A3(\b_l[6] ),
    .A4(\b_l[7] ),
    .B1(_09330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09336_));
 sky130_fd_sc_hd__and4_2 _18475_ (.A(_09334_),
    .B(_09335_),
    .C(\a_l[3] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09337_));
 sky130_fd_sc_hd__a22o_2 _18476_ (.A1(\a_l[3] ),
    .A2(\b_l[8] ),
    .B1(_09334_),
    .B2(_09335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09338_));
 sky130_fd_sc_hd__o221ai_2 _18477_ (.A1(_09188_),
    .A2(_09264_),
    .B1(_04260_),
    .B2(_06605_),
    .C1(_09334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09339_));
 sky130_fd_sc_hd__a21o_2 _18478_ (.A1(_09334_),
    .A2(_09335_),
    .B1(_09330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09341_));
 sky130_fd_sc_hd__nand2_2 _18479_ (.A(_09338_),
    .B(_09327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09342_));
 sky130_fd_sc_hd__o211ai_2 _18480_ (.A1(_09333_),
    .A2(_09336_),
    .B1(_09327_),
    .C1(_09338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09343_));
 sky130_fd_sc_hd__nand3_2 _18481_ (.A(_09328_),
    .B(_09339_),
    .C(_09341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09344_));
 sky130_fd_sc_hd__a32o_2 _18482_ (.A1(\a_l[3] ),
    .A2(\a_l[4] ),
    .A3(_04259_),
    .B1(_09269_),
    .B2(_09274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09345_));
 sky130_fd_sc_hd__a21boi_2 _18483_ (.A1(_09343_),
    .A2(_09344_),
    .B1_N(_09345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09346_));
 sky130_fd_sc_hd__o2111a_2 _18484_ (.A1(_09270_),
    .A2(_09273_),
    .B1(_09276_),
    .C1(_09343_),
    .D1(_09344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09347_));
 sky130_fd_sc_hd__a21o_2 _18485_ (.A1(_09343_),
    .A2(_09344_),
    .B1(_09345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09348_));
 sky130_fd_sc_hd__o211ai_2 _18486_ (.A1(_09337_),
    .A2(_09342_),
    .B1(_09344_),
    .C1(_09345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09349_));
 sky130_fd_sc_hd__nand2_2 _18487_ (.A(_09348_),
    .B(_09349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09350_));
 sky130_fd_sc_hd__a32oi_2 _18488_ (.A1(_09233_),
    .A2(_09240_),
    .A3(_09241_),
    .B1(_09254_),
    .B2(_09256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09352_));
 sky130_fd_sc_hd__a32oi_2 _18489_ (.A1(_09232_),
    .A2(_09244_),
    .A3(_09245_),
    .B1(_09259_),
    .B2(_09243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09353_));
 sky130_fd_sc_hd__nand2_2 _18490_ (.A(\b_l[5] ),
    .B(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_2 _18491_ (.A(\b_l[3] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09355_));
 sky130_fd_sc_hd__nand2_2 _18492_ (.A(\b_l[4] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_2 _18493_ (.A(_09355_),
    .B(_09356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09357_));
 sky130_fd_sc_hd__nand2_2 _18494_ (.A(\b_l[4] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09358_));
 sky130_fd_sc_hd__and4_2 _18495_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[7] ),
    .D(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09359_));
 sky130_fd_sc_hd__nand4_2 _18496_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[7] ),
    .D(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09360_));
 sky130_fd_sc_hd__a22oi_2 _18497_ (.A1(\b_l[5] ),
    .A2(\a_l[6] ),
    .B1(_09357_),
    .B2(_09360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09361_));
 sky130_fd_sc_hd__o21ba_2 _18498_ (.A1(_04182_),
    .A2(_06867_),
    .B1_N(_09354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09363_));
 sky130_fd_sc_hd__a21o_2 _18499_ (.A1(_09363_),
    .A2(_09357_),
    .B1(_09361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09364_));
 sky130_fd_sc_hd__a21oi_2 _18500_ (.A1(_09363_),
    .A2(_09357_),
    .B1(_09361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09365_));
 sky130_fd_sc_hd__o21a_2 _18501_ (.A1(_04134_),
    .A2(_07100_),
    .B1(_09234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09366_));
 sky130_fd_sc_hd__o21ai_2 _18502_ (.A1(_04134_),
    .A2(_07100_),
    .B1(_09234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09367_));
 sky130_fd_sc_hd__a21oi_2 _18503_ (.A1(_09234_),
    .A2(_09239_),
    .B1(_09237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09368_));
 sky130_fd_sc_hd__nand2_2 _18504_ (.A(\b_l[2] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09369_));
 sky130_fd_sc_hd__nand2_2 _18505_ (.A(\b_l[1] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09370_));
 sky130_fd_sc_hd__nand2_2 _18506_ (.A(\b_l[0] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09371_));
 sky130_fd_sc_hd__a22oi_2 _18507_ (.A1(\b_l[1] ),
    .A2(\a_l[10] ),
    .B1(\a_l[11] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09372_));
 sky130_fd_sc_hd__nand2_2 _18508_ (.A(_09370_),
    .B(_09371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09374_));
 sky130_fd_sc_hd__nand4_2 _18509_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[10] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09375_));
 sky130_fd_sc_hd__o221ai_2 _18510_ (.A1(_09155_),
    .A2(_09275_),
    .B1(_04134_),
    .B2(_07234_),
    .C1(_09374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09376_));
 sky130_fd_sc_hd__a21o_2 _18511_ (.A1(_09374_),
    .A2(_09375_),
    .B1(_09369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09377_));
 sky130_fd_sc_hd__o2bb2ai_2 _18512_ (.A1_N(_09374_),
    .A2_N(_09375_),
    .B1(_09155_),
    .B2(_09275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09378_));
 sky130_fd_sc_hd__nand3_2 _18513_ (.A(_09375_),
    .B(\a_l[9] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09379_));
 sky130_fd_sc_hd__o211ai_2 _18514_ (.A1(_09237_),
    .A2(_09366_),
    .B1(_09376_),
    .C1(_09377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09380_));
 sky130_fd_sc_hd__o211ai_2 _18515_ (.A1(_09379_),
    .A2(_09372_),
    .B1(_09367_),
    .C1(_09378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09381_));
 sky130_fd_sc_hd__o211ai_2 _18516_ (.A1(_09379_),
    .A2(_09372_),
    .B1(_09368_),
    .C1(_09378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09382_));
 sky130_fd_sc_hd__nand3_2 _18517_ (.A(_09365_),
    .B(_09380_),
    .C(_09382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09383_));
 sky130_fd_sc_hd__a21o_2 _18518_ (.A1(_09380_),
    .A2(_09382_),
    .B1(_09365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09385_));
 sky130_fd_sc_hd__nand3_2 _18519_ (.A(_09385_),
    .B(_09353_),
    .C(_09383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09386_));
 sky130_fd_sc_hd__inv_2 _18520_ (.A(_09386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09387_));
 sky130_fd_sc_hd__and3_2 _18521_ (.A(_09364_),
    .B(_09380_),
    .C(_09382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09388_));
 sky130_fd_sc_hd__o211ai_2 _18522_ (.A1(_09237_),
    .A2(_09381_),
    .B1(_09380_),
    .C1(_09364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09389_));
 sky130_fd_sc_hd__a21o_2 _18523_ (.A1(_09380_),
    .A2(_09382_),
    .B1(_09364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09390_));
 sky130_fd_sc_hd__o21ai_2 _18524_ (.A1(_09246_),
    .A2(_09352_),
    .B1(_09390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09391_));
 sky130_fd_sc_hd__a2bb2oi_2 _18525_ (.A1_N(_09246_),
    .A2_N(_09352_),
    .B1(_09383_),
    .B2(_09385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09392_));
 sky130_fd_sc_hd__o211ai_2 _18526_ (.A1(_09246_),
    .A2(_09352_),
    .B1(_09389_),
    .C1(_09390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09393_));
 sky130_fd_sc_hd__nand2_2 _18527_ (.A(_09386_),
    .B(_09393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09394_));
 sky130_fd_sc_hd__nand2_2 _18528_ (.A(_09393_),
    .B(_09350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09396_));
 sky130_fd_sc_hd__o211ai_2 _18529_ (.A1(_09388_),
    .A2(_09391_),
    .B1(_09350_),
    .C1(_09386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09397_));
 sky130_fd_sc_hd__o21ai_2 _18530_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09398_));
 sky130_fd_sc_hd__nand2_2 _18531_ (.A(_09394_),
    .B(_09350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09399_));
 sky130_fd_sc_hd__o211ai_2 _18532_ (.A1(_09346_),
    .A2(_09347_),
    .B1(_09386_),
    .C1(_09393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09400_));
 sky130_fd_sc_hd__o211a_2 _18533_ (.A1(_09396_),
    .A2(_09387_),
    .B1(_09326_),
    .C1(_09398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09401_));
 sky130_fd_sc_hd__o211ai_2 _18534_ (.A1(_09396_),
    .A2(_09387_),
    .B1(_09326_),
    .C1(_09398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09402_));
 sky130_fd_sc_hd__nand3_2 _18535_ (.A(_09399_),
    .B(_09400_),
    .C(_09325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09403_));
 sky130_fd_sc_hd__nand2_2 _18536_ (.A(\a_l[2] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09404_));
 sky130_fd_sc_hd__nand4_2 _18537_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09405_));
 sky130_fd_sc_hd__a22oi_2 _18538_ (.A1(\a_l[2] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09407_));
 sky130_fd_sc_hd__nand2_2 _18539_ (.A(_09216_),
    .B(_09404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_2 _18540_ (.A(\a_l[0] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09409_));
 sky130_fd_sc_hd__a21oi_2 _18541_ (.A1(_09405_),
    .A2(_09408_),
    .B1(_09409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09410_));
 sky130_fd_sc_hd__o221a_2 _18542_ (.A1(_09166_),
    .A2(_09308_),
    .B1(_04555_),
    .B2(_06441_),
    .C1(_09408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09411_));
 sky130_fd_sc_hd__o2111ai_2 _18543_ (.A1(_09410_),
    .A2(_09411_),
    .B1(\b_l[9] ),
    .C1(\b_l[10] ),
    .D1(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09412_));
 sky130_fd_sc_hd__a211o_2 _18544_ (.A1(\b_l[10] ),
    .A2(_09217_),
    .B1(_09410_),
    .C1(_09411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09413_));
 sky130_fd_sc_hd__nand2_2 _18545_ (.A(_09412_),
    .B(_09413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09414_));
 sky130_fd_sc_hd__a31o_2 _18546_ (.A1(_09118_),
    .A2(_09123_),
    .A3(_09283_),
    .B1(_09281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09415_));
 sky130_fd_sc_hd__nor2_2 _18547_ (.A(_09414_),
    .B(_09415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09416_));
 sky130_fd_sc_hd__nand2_2 _18548_ (.A(_09414_),
    .B(_09415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09418_));
 sky130_fd_sc_hd__a21oi_2 _18549_ (.A1(_09412_),
    .A2(_09413_),
    .B1(_09415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09419_));
 sky130_fd_sc_hd__and3_2 _18550_ (.A(_09412_),
    .B(_09413_),
    .C(_09415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09420_));
 sky130_fd_sc_hd__and2b_2 _18551_ (.A_N(_09416_),
    .B(_09418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09421_));
 sky130_fd_sc_hd__nor2_2 _18552_ (.A(_09419_),
    .B(_09420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09422_));
 sky130_fd_sc_hd__a21oi_2 _18553_ (.A1(_09402_),
    .A2(_09403_),
    .B1(_09421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09423_));
 sky130_fd_sc_hd__a21o_2 _18554_ (.A1(_09402_),
    .A2(_09403_),
    .B1(_09421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09424_));
 sky130_fd_sc_hd__o211ai_2 _18555_ (.A1(_09419_),
    .A2(_09420_),
    .B1(_09402_),
    .C1(_09403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09425_));
 sky130_fd_sc_hd__o2bb2ai_2 _18556_ (.A1_N(_09402_),
    .A2_N(_09403_),
    .B1(_09419_),
    .B2(_09420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09426_));
 sky130_fd_sc_hd__nand3_2 _18557_ (.A(_09402_),
    .B(_09403_),
    .C(_09422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_2 _18558_ (.A(_09323_),
    .B(_09425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09429_));
 sky130_fd_sc_hd__nand3_2 _18559_ (.A(_09424_),
    .B(_09425_),
    .C(_09323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09430_));
 sky130_fd_sc_hd__nand3_2 _18560_ (.A(_09324_),
    .B(_09426_),
    .C(_09427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09431_));
 sky130_fd_sc_hd__o2bb2ai_2 _18561_ (.A1_N(_09430_),
    .A2_N(_09431_),
    .B1(_09219_),
    .B2(_09222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09432_));
 sky130_fd_sc_hd__nand2_2 _18562_ (.A(_09431_),
    .B(_09223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09433_));
 sky130_fd_sc_hd__o211ai_2 _18563_ (.A1(_09423_),
    .A2(_09429_),
    .B1(_09223_),
    .C1(_09431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09434_));
 sky130_fd_sc_hd__a22oi_2 _18564_ (.A1(_09303_),
    .A2(_09299_),
    .B1(_09191_),
    .B2(_09306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09435_));
 sky130_fd_sc_hd__a21o_2 _18565_ (.A1(_09432_),
    .A2(_09434_),
    .B1(_09435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09436_));
 sky130_fd_sc_hd__nand3_2 _18566_ (.A(_09432_),
    .B(_09434_),
    .C(_09435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09437_));
 sky130_fd_sc_hd__and2_2 _18567_ (.A(_09436_),
    .B(_09437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09438_));
 sky130_fd_sc_hd__a21oi_2 _18568_ (.A1(_09436_),
    .A2(_09437_),
    .B1(_09313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09440_));
 sky130_fd_sc_hd__a21o_2 _18569_ (.A1(_09313_),
    .A2(_09436_),
    .B1(_09440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09441_));
 sky130_fd_sc_hd__nand2_2 _18570_ (.A(_09322_),
    .B(_09441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09442_));
 sky130_fd_sc_hd__o211a_2 _18571_ (.A1(_09322_),
    .A2(_09440_),
    .B1(_09442_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00381_));
 sky130_fd_sc_hd__o2bb2ai_2 _18572_ (.A1_N(_09223_),
    .A2_N(_09431_),
    .B1(_09429_),
    .B2(_09423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09443_));
 sky130_fd_sc_hd__a21boi_2 _18573_ (.A1(_09223_),
    .A2(_09431_),
    .B1_N(_09430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09444_));
 sky130_fd_sc_hd__o2bb2ai_2 _18574_ (.A1_N(_09350_),
    .A2_N(_09386_),
    .B1(_09388_),
    .B2(_09391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09445_));
 sky130_fd_sc_hd__a21oi_2 _18575_ (.A1(_09386_),
    .A2(_09350_),
    .B1(_09392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09446_));
 sky130_fd_sc_hd__o21ai_2 _18576_ (.A1(_04182_),
    .A2(_06867_),
    .B1(_09354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09447_));
 sky130_fd_sc_hd__a21oi_2 _18577_ (.A1(_09355_),
    .A2(_09356_),
    .B1(_09354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09448_));
 sky130_fd_sc_hd__nand2_2 _18578_ (.A(_09357_),
    .B(_09447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09450_));
 sky130_fd_sc_hd__and2_2 _18579_ (.A(\a_l[4] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09451_));
 sky130_fd_sc_hd__nand2_2 _18580_ (.A(\a_l[5] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09452_));
 sky130_fd_sc_hd__nand2_2 _18581_ (.A(\a_l[6] ),
    .B(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09453_));
 sky130_fd_sc_hd__a22o_2 _18582_ (.A1(\a_l[6] ),
    .A2(\b_l[6] ),
    .B1(\b_l[7] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09454_));
 sky130_fd_sc_hd__nand3_2 _18583_ (.A(_09453_),
    .B(\b_l[7] ),
    .C(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09455_));
 sky130_fd_sc_hd__nand3_2 _18584_ (.A(_09452_),
    .B(\b_l[6] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09456_));
 sky130_fd_sc_hd__o221ai_2 _18585_ (.A1(_09199_),
    .A2(_09264_),
    .B1(_04260_),
    .B2(_06681_),
    .C1(_09454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09457_));
 sky130_fd_sc_hd__nand4_2 _18586_ (.A(_09455_),
    .B(_09456_),
    .C(\a_l[4] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09458_));
 sky130_fd_sc_hd__o211ai_2 _18587_ (.A1(_09199_),
    .A2(_09264_),
    .B1(_09455_),
    .C1(_09456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09459_));
 sky130_fd_sc_hd__o211ai_2 _18588_ (.A1(_04260_),
    .A2(_06681_),
    .B1(_09451_),
    .C1(_09454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09461_));
 sky130_fd_sc_hd__o211ai_2 _18589_ (.A1(_09359_),
    .A2(_09448_),
    .B1(_09459_),
    .C1(_09461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09462_));
 sky130_fd_sc_hd__and3_2 _18590_ (.A(_09450_),
    .B(_09457_),
    .C(_09458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09463_));
 sky130_fd_sc_hd__nand3_2 _18591_ (.A(_09450_),
    .B(_09457_),
    .C(_09458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09464_));
 sky130_fd_sc_hd__o32a_2 _18592_ (.A1(_09199_),
    .A2(_09210_),
    .A3(_04260_),
    .B1(_09264_),
    .B2(_09188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09465_));
 sky130_fd_sc_hd__a32o_2 _18593_ (.A1(\a_l[4] ),
    .A2(\a_l[5] ),
    .A3(_04259_),
    .B1(\b_l[8] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09466_));
 sky130_fd_sc_hd__o32a_2 _18594_ (.A1(_09199_),
    .A2(_09210_),
    .A3(_04260_),
    .B1(_09330_),
    .B2(_09333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09467_));
 sky130_fd_sc_hd__and3_2 _18595_ (.A(_09462_),
    .B(_09464_),
    .C(_09467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09468_));
 sky130_fd_sc_hd__a21oi_2 _18596_ (.A1(_09462_),
    .A2(_09464_),
    .B1(_09467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09469_));
 sky130_fd_sc_hd__o2bb2ai_2 _18597_ (.A1_N(_09462_),
    .A2_N(_09464_),
    .B1(_09465_),
    .B2(_09333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09470_));
 sky130_fd_sc_hd__nand4_2 _18598_ (.A(_09334_),
    .B(_09462_),
    .C(_09464_),
    .D(_09466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09472_));
 sky130_fd_sc_hd__nand2_2 _18599_ (.A(_09470_),
    .B(_09472_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09473_));
 sky130_fd_sc_hd__o2bb2ai_2 _18600_ (.A1_N(_09365_),
    .A2_N(_09380_),
    .B1(_09381_),
    .B2(_09237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09474_));
 sky130_fd_sc_hd__a21boi_2 _18601_ (.A1(_09365_),
    .A2(_09380_),
    .B1_N(_09382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09475_));
 sky130_fd_sc_hd__o21a_2 _18602_ (.A1(_04134_),
    .A2(_07234_),
    .B1(_09369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09476_));
 sky130_fd_sc_hd__o21ai_2 _18603_ (.A1(_09369_),
    .A2(_09372_),
    .B1(_09375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09477_));
 sky130_fd_sc_hd__nand2_2 _18604_ (.A(\b_l[1] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09478_));
 sky130_fd_sc_hd__nand2_2 _18605_ (.A(\b_l[0] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_2 _18606_ (.A(_09478_),
    .B(_09479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09480_));
 sky130_fd_sc_hd__nand2_2 _18607_ (.A(\b_l[1] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09481_));
 sky130_fd_sc_hd__and4_2 _18608_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[11] ),
    .D(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09483_));
 sky130_fd_sc_hd__nand4_2 _18609_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[11] ),
    .D(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09484_));
 sky130_fd_sc_hd__nand2_2 _18610_ (.A(_09480_),
    .B(_09484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09485_));
 sky130_fd_sc_hd__nor2_2 _18611_ (.A(_09155_),
    .B(_09286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09486_));
 sky130_fd_sc_hd__nand2_2 _18612_ (.A(\b_l[2] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09487_));
 sky130_fd_sc_hd__a22o_2 _18613_ (.A1(\b_l[2] ),
    .A2(\a_l[10] ),
    .B1(_09480_),
    .B2(_09484_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09488_));
 sky130_fd_sc_hd__o311a_2 _18614_ (.A1(_09297_),
    .A2(_09319_),
    .A3(_04134_),
    .B1(_09480_),
    .C1(_09486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09489_));
 sky130_fd_sc_hd__o2111ai_2 _18615_ (.A1(_09371_),
    .A2(_09481_),
    .B1(\b_l[2] ),
    .C1(\a_l[10] ),
    .D1(_09480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09490_));
 sky130_fd_sc_hd__o221ai_2 _18616_ (.A1(_09155_),
    .A2(_09286_),
    .B1(_09371_),
    .B2(_09481_),
    .C1(_09480_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09491_));
 sky130_fd_sc_hd__nand2_2 _18617_ (.A(_09485_),
    .B(_09486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09492_));
 sky130_fd_sc_hd__o211ai_2 _18618_ (.A1(_09372_),
    .A2(_09476_),
    .B1(_09491_),
    .C1(_09492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_2 _18619_ (.A(_09488_),
    .B(_09477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09495_));
 sky130_fd_sc_hd__nand3_2 _18620_ (.A(_09488_),
    .B(_09490_),
    .C(_09477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09496_));
 sky130_fd_sc_hd__and2_2 _18621_ (.A(\b_l[5] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09497_));
 sky130_fd_sc_hd__nand2_2 _18622_ (.A(\b_l[5] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_2 _18623_ (.A(\b_l[3] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09499_));
 sky130_fd_sc_hd__a22oi_2 _18624_ (.A1(\b_l[4] ),
    .A2(\a_l[8] ),
    .B1(\a_l[9] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_2 _18625_ (.A(_09358_),
    .B(_09499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09501_));
 sky130_fd_sc_hd__nand4_2 _18626_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[8] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09502_));
 sky130_fd_sc_hd__o221a_2 _18627_ (.A1(_09220_),
    .A2(_09242_),
    .B1(_04182_),
    .B2(_06985_),
    .C1(_09501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09503_));
 sky130_fd_sc_hd__a21oi_2 _18628_ (.A1(_09501_),
    .A2(_09502_),
    .B1(_09498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09505_));
 sky130_fd_sc_hd__a21oi_2 _18629_ (.A1(_09501_),
    .A2(_09502_),
    .B1(_09497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09506_));
 sky130_fd_sc_hd__and3_2 _18630_ (.A(_09501_),
    .B(_09502_),
    .C(_09497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09507_));
 sky130_fd_sc_hd__nor2_2 _18631_ (.A(_09506_),
    .B(_09507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09508_));
 sky130_fd_sc_hd__o211ai_2 _18632_ (.A1(_09503_),
    .A2(_09505_),
    .B1(_09494_),
    .C1(_09496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09509_));
 sky130_fd_sc_hd__o2bb2ai_2 _18633_ (.A1_N(_09494_),
    .A2_N(_09496_),
    .B1(_09506_),
    .B2(_09507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09510_));
 sky130_fd_sc_hd__and3_2 _18634_ (.A(_09510_),
    .B(_09474_),
    .C(_09509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09511_));
 sky130_fd_sc_hd__nand3_2 _18635_ (.A(_09510_),
    .B(_09474_),
    .C(_09509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09512_));
 sky130_fd_sc_hd__o211ai_2 _18636_ (.A1(_09506_),
    .A2(_09507_),
    .B1(_09494_),
    .C1(_09496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09513_));
 sky130_fd_sc_hd__inv_2 _18637_ (.A(_09513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09514_));
 sky130_fd_sc_hd__o2bb2ai_2 _18638_ (.A1_N(_09494_),
    .A2_N(_09496_),
    .B1(_09503_),
    .B2(_09505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09516_));
 sky130_fd_sc_hd__nand2_2 _18639_ (.A(_09475_),
    .B(_09516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09517_));
 sky130_fd_sc_hd__nand3_2 _18640_ (.A(_09475_),
    .B(_09513_),
    .C(_09516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09518_));
 sky130_fd_sc_hd__nand2_2 _18641_ (.A(_09512_),
    .B(_09518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09519_));
 sky130_fd_sc_hd__a31oi_2 _18642_ (.A1(_09475_),
    .A2(_09513_),
    .A3(_09516_),
    .B1(_09473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09520_));
 sky130_fd_sc_hd__o21ai_2 _18643_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09521_));
 sky130_fd_sc_hd__o211a_2 _18644_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09512_),
    .C1(_09518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09522_));
 sky130_fd_sc_hd__nand2_2 _18645_ (.A(_09519_),
    .B(_09473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09523_));
 sky130_fd_sc_hd__o21ai_2 _18646_ (.A1(_09468_),
    .A2(_09469_),
    .B1(_09519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09524_));
 sky130_fd_sc_hd__o211ai_2 _18647_ (.A1(_09514_),
    .A2(_09517_),
    .B1(_09473_),
    .C1(_09512_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_2 _18648_ (.A(_09446_),
    .B(_09523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09527_));
 sky130_fd_sc_hd__a21oi_2 _18649_ (.A1(_09524_),
    .A2(_09525_),
    .B1(_09445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09528_));
 sky130_fd_sc_hd__o211ai_2 _18650_ (.A1(_09521_),
    .A2(_09511_),
    .B1(_09446_),
    .C1(_09523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09529_));
 sky130_fd_sc_hd__nand3_2 _18651_ (.A(_09524_),
    .B(_09525_),
    .C(_09445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_2 _18652_ (.A1(_09405_),
    .A2(_09409_),
    .B1(_09407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09531_));
 sky130_fd_sc_hd__a21o_2 _18653_ (.A1(_09405_),
    .A2(_09409_),
    .B1(_09407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09532_));
 sky130_fd_sc_hd__nand2_2 _18654_ (.A(\a_l[1] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_2 _18655_ (.A(\a_l[2] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09534_));
 sky130_fd_sc_hd__nand2_2 _18656_ (.A(\a_l[3] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09535_));
 sky130_fd_sc_hd__a22oi_2 _18657_ (.A1(\a_l[3] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_2 _18658_ (.A(_09534_),
    .B(_09535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09538_));
 sky130_fd_sc_hd__nand4_2 _18659_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09539_));
 sky130_fd_sc_hd__a22o_2 _18660_ (.A1(\a_l[1] ),
    .A2(\b_l[11] ),
    .B1(_09538_),
    .B2(_09539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09540_));
 sky130_fd_sc_hd__nand4_2 _18661_ (.A(_09538_),
    .B(_09539_),
    .C(\a_l[1] ),
    .D(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09541_));
 sky130_fd_sc_hd__a21o_2 _18662_ (.A1(_09538_),
    .A2(_09539_),
    .B1(_09533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09542_));
 sky130_fd_sc_hd__nand3_2 _18663_ (.A(_09533_),
    .B(_09538_),
    .C(_09539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09543_));
 sky130_fd_sc_hd__nand3_2 _18664_ (.A(_09532_),
    .B(_09542_),
    .C(_09543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09544_));
 sky130_fd_sc_hd__and3_2 _18665_ (.A(_09540_),
    .B(_09541_),
    .C(_09531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09545_));
 sky130_fd_sc_hd__nand3_2 _18666_ (.A(_09540_),
    .B(_09541_),
    .C(_09531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09546_));
 sky130_fd_sc_hd__o2bb2ai_2 _18667_ (.A1_N(_09544_),
    .A2_N(_09546_),
    .B1(_09166_),
    .B2(_09329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09547_));
 sky130_fd_sc_hd__nand3_2 _18668_ (.A(_09544_),
    .B(\b_l[12] ),
    .C(\a_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09549_));
 sky130_fd_sc_hd__nand4_2 _18669_ (.A(_09544_),
    .B(_09546_),
    .C(\a_l[0] ),
    .D(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09550_));
 sky130_fd_sc_hd__o2bb2ai_2 _18670_ (.A1_N(_09345_),
    .A2_N(_09344_),
    .B1(_09342_),
    .B2(_09337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09551_));
 sky130_fd_sc_hd__a21oi_2 _18671_ (.A1(_09547_),
    .A2(_09550_),
    .B1(_09551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09552_));
 sky130_fd_sc_hd__a21o_2 _18672_ (.A1(_09547_),
    .A2(_09550_),
    .B1(_09551_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09553_));
 sky130_fd_sc_hd__o211a_2 _18673_ (.A1(_09545_),
    .A2(_09549_),
    .B1(_09551_),
    .C1(_09547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09554_));
 sky130_fd_sc_hd__o211ai_2 _18674_ (.A1(_09545_),
    .A2(_09549_),
    .B1(_09551_),
    .C1(_09547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09555_));
 sky130_fd_sc_hd__o2111a_2 _18675_ (.A1(_09410_),
    .A2(_09411_),
    .B1(\b_l[10] ),
    .C1(_09217_),
    .D1(_09553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09556_));
 sky130_fd_sc_hd__a21oi_2 _18676_ (.A1(_09553_),
    .A2(_09555_),
    .B1(_09412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09557_));
 sky130_fd_sc_hd__o21bai_2 _18677_ (.A1(_09552_),
    .A2(_09554_),
    .B1_N(_09412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09558_));
 sky130_fd_sc_hd__and3_2 _18678_ (.A(_09412_),
    .B(_09553_),
    .C(_09555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09560_));
 sky130_fd_sc_hd__nand3_2 _18679_ (.A(_09412_),
    .B(_09553_),
    .C(_09555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09561_));
 sky130_fd_sc_hd__nand2_2 _18680_ (.A(_09558_),
    .B(_09561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09562_));
 sky130_fd_sc_hd__o2bb2ai_2 _18681_ (.A1_N(_09529_),
    .A2_N(_09530_),
    .B1(_09557_),
    .B2(_09560_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09563_));
 sky130_fd_sc_hd__nand4_2 _18682_ (.A(_09529_),
    .B(_09530_),
    .C(_09558_),
    .D(_09561_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09564_));
 sky130_fd_sc_hd__a21oi_2 _18683_ (.A1(_09529_),
    .A2(_09530_),
    .B1(_09562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09565_));
 sky130_fd_sc_hd__a21o_2 _18684_ (.A1(_09529_),
    .A2(_09530_),
    .B1(_09562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09566_));
 sky130_fd_sc_hd__nand3_2 _18685_ (.A(_09529_),
    .B(_09530_),
    .C(_09562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09567_));
 sky130_fd_sc_hd__a31oi_2 _18686_ (.A1(_09399_),
    .A2(_09400_),
    .A3(_09325_),
    .B1(_09421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09568_));
 sky130_fd_sc_hd__nand2_2 _18687_ (.A(_09403_),
    .B(_09422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09569_));
 sky130_fd_sc_hd__a32oi_2 _18688_ (.A1(_09326_),
    .A2(_09397_),
    .A3(_09398_),
    .B1(_09403_),
    .B2(_09422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09571_));
 sky130_fd_sc_hd__o211ai_2 _18689_ (.A1(_09401_),
    .A2(_09568_),
    .B1(_09564_),
    .C1(_09563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09572_));
 sky130_fd_sc_hd__nand3_2 _18690_ (.A(_09402_),
    .B(_09567_),
    .C(_09569_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09573_));
 sky130_fd_sc_hd__nand3_2 _18691_ (.A(_09566_),
    .B(_09571_),
    .C(_09567_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09574_));
 sky130_fd_sc_hd__o21ai_2 _18692_ (.A1(_09565_),
    .A2(_09573_),
    .B1(_09572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09575_));
 sky130_fd_sc_hd__o211ai_2 _18693_ (.A1(_09565_),
    .A2(_09573_),
    .B1(_09572_),
    .C1(_09416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09576_));
 sky130_fd_sc_hd__o2bb2ai_2 _18694_ (.A1_N(_09572_),
    .A2_N(_09574_),
    .B1(_09414_),
    .B2(_09415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09577_));
 sky130_fd_sc_hd__o221ai_2 _18695_ (.A1(_09414_),
    .A2(_09415_),
    .B1(_09565_),
    .B2(_09573_),
    .C1(_09572_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09578_));
 sky130_fd_sc_hd__nand2_2 _18696_ (.A(_09575_),
    .B(_09416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09579_));
 sky130_fd_sc_hd__nand3_2 _18697_ (.A(_09444_),
    .B(_09578_),
    .C(_09579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09580_));
 sky130_fd_sc_hd__a22oi_2 _18698_ (.A1(_09430_),
    .A2(_09433_),
    .B1(_09578_),
    .B2(_09579_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09582_));
 sky130_fd_sc_hd__nand3_2 _18699_ (.A(_09443_),
    .B(_09576_),
    .C(_09577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09583_));
 sky130_fd_sc_hd__nand2_2 _18700_ (.A(_09580_),
    .B(_09583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09584_));
 sky130_fd_sc_hd__a21boi_2 _18701_ (.A1(_09580_),
    .A2(_09583_),
    .B1_N(_09437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09585_));
 sky130_fd_sc_hd__a31oi_2 _18702_ (.A1(_09443_),
    .A2(_09576_),
    .A3(_09577_),
    .B1(_09437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09586_));
 sky130_fd_sc_hd__a21oi_2 _18703_ (.A1(_09586_),
    .A2(_09580_),
    .B1(_09585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09587_));
 sky130_fd_sc_hd__a21o_2 _18704_ (.A1(_09586_),
    .A2(_09580_),
    .B1(_09585_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09588_));
 sky130_fd_sc_hd__a22oi_2 _18705_ (.A1(_09207_),
    .A2(_09312_),
    .B1(_09436_),
    .B2(_09313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09589_));
 sky130_fd_sc_hd__o21ai_2 _18706_ (.A1(_09315_),
    .A2(_09320_),
    .B1(_09589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09590_));
 sky130_fd_sc_hd__o2bb2a_2 _18707_ (.A1_N(_09313_),
    .A2_N(_09436_),
    .B1(_09440_),
    .B2(_09322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09591_));
 sky130_fd_sc_hd__o21a_2 _18708_ (.A1(_09588_),
    .A2(_09591_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09593_));
 sky130_fd_sc_hd__a21boi_2 _18709_ (.A1(_09588_),
    .A2(_09591_),
    .B1_N(_09593_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00382_));
 sky130_fd_sc_hd__o21a_2 _18710_ (.A1(_09333_),
    .A2(_09465_),
    .B1(_09462_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09594_));
 sky130_fd_sc_hd__a21oi_2 _18711_ (.A1(_09462_),
    .A2(_09467_),
    .B1(_09463_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09595_));
 sky130_fd_sc_hd__and3_2 _18712_ (.A(\a_l[1] ),
    .B(\a_l[0] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09596_));
 sky130_fd_sc_hd__o2bb2a_2 _18713_ (.A1_N(\a_l[1] ),
    .A2_N(\b_l[12] ),
    .B1(_09351_),
    .B2(_09166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09597_));
 sky130_fd_sc_hd__a21oi_2 _18714_ (.A1(_05043_),
    .A2(_06401_),
    .B1(_09597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09598_));
 sky130_fd_sc_hd__o21ai_2 _18715_ (.A1(_09534_),
    .A2(_09535_),
    .B1(_09533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09599_));
 sky130_fd_sc_hd__o21ai_2 _18716_ (.A1(_09533_),
    .A2(_09536_),
    .B1(_09539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09600_));
 sky130_fd_sc_hd__o21a_2 _18717_ (.A1(_09533_),
    .A2(_09536_),
    .B1(_09539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09601_));
 sky130_fd_sc_hd__nand2_2 _18718_ (.A(\a_l[3] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09603_));
 sky130_fd_sc_hd__nand2_2 _18719_ (.A(\a_l[4] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09604_));
 sky130_fd_sc_hd__a22oi_2 _18720_ (.A1(\a_l[4] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09605_));
 sky130_fd_sc_hd__nand2_2 _18721_ (.A(_09603_),
    .B(_09604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09606_));
 sky130_fd_sc_hd__nor2_2 _18722_ (.A(_04555_),
    .B(_06521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09607_));
 sky130_fd_sc_hd__nand4_2 _18723_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09608_));
 sky130_fd_sc_hd__nand2_2 _18724_ (.A(\a_l[2] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09609_));
 sky130_fd_sc_hd__o21ai_2 _18725_ (.A1(_09605_),
    .A2(_09607_),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09610_));
 sky130_fd_sc_hd__a41o_2 _18726_ (.A1(\a_l[3] ),
    .A2(\a_l[4] ),
    .A3(\b_l[9] ),
    .A4(\b_l[10] ),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09611_));
 sky130_fd_sc_hd__o211ai_2 _18727_ (.A1(_09605_),
    .A2(_09611_),
    .B1(_09600_),
    .C1(_09610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09612_));
 sky130_fd_sc_hd__a21oi_2 _18728_ (.A1(_09606_),
    .A2(_09608_),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09614_));
 sky130_fd_sc_hd__a21o_2 _18729_ (.A1(_09606_),
    .A2(_09608_),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09615_));
 sky130_fd_sc_hd__o22a_2 _18730_ (.A1(_09144_),
    .A2(_09308_),
    .B1(_04555_),
    .B2(_06521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09616_));
 sky130_fd_sc_hd__o21ai_2 _18731_ (.A1(_04555_),
    .A2(_06521_),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09617_));
 sky130_fd_sc_hd__o2bb2ai_2 _18732_ (.A1_N(_09538_),
    .A2_N(_09599_),
    .B1(_09605_),
    .B2(_09617_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09618_));
 sky130_fd_sc_hd__o211ai_2 _18733_ (.A1(_09617_),
    .A2(_09605_),
    .B1(_09601_),
    .C1(_09615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09619_));
 sky130_fd_sc_hd__o211a_2 _18734_ (.A1(_09614_),
    .A2(_09618_),
    .B1(_09598_),
    .C1(_09612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09620_));
 sky130_fd_sc_hd__o211ai_2 _18735_ (.A1(_09614_),
    .A2(_09618_),
    .B1(_09598_),
    .C1(_09612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09621_));
 sky130_fd_sc_hd__a21oi_2 _18736_ (.A1(_09612_),
    .A2(_09619_),
    .B1(_09598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09622_));
 sky130_fd_sc_hd__a2bb2o_2 _18737_ (.A1_N(_09596_),
    .A2_N(_09597_),
    .B1(_09612_),
    .B2(_09619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09623_));
 sky130_fd_sc_hd__and3_2 _18738_ (.A(_09595_),
    .B(_09621_),
    .C(_09623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09625_));
 sky130_fd_sc_hd__nand3_2 _18739_ (.A(_09595_),
    .B(_09621_),
    .C(_09623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09626_));
 sky130_fd_sc_hd__o22ai_2 _18740_ (.A1(_09463_),
    .A2(_09594_),
    .B1(_09620_),
    .B2(_09622_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09627_));
 sky130_fd_sc_hd__a31o_2 _18741_ (.A1(\a_l[0] ),
    .A2(\b_l[12] ),
    .A3(_09544_),
    .B1(_09545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09628_));
 sky130_fd_sc_hd__and3_2 _18742_ (.A(_09626_),
    .B(_09627_),
    .C(_09628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09629_));
 sky130_fd_sc_hd__nand3_2 _18743_ (.A(_09626_),
    .B(_09627_),
    .C(_09628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09630_));
 sky130_fd_sc_hd__a21o_2 _18744_ (.A1(_09626_),
    .A2(_09627_),
    .B1(_09628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09631_));
 sky130_fd_sc_hd__a22o_2 _18745_ (.A1(_09546_),
    .A2(_09549_),
    .B1(_09626_),
    .B2(_09627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09632_));
 sky130_fd_sc_hd__nand4_2 _18746_ (.A(_09546_),
    .B(_09549_),
    .C(_09626_),
    .D(_09627_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_2 _18747_ (.A(_09632_),
    .B(_09633_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09634_));
 sky130_fd_sc_hd__o2bb2ai_2 _18748_ (.A1_N(_09473_),
    .A2_N(_09512_),
    .B1(_09514_),
    .B2(_09517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09636_));
 sky130_fd_sc_hd__o2bb2ai_2 _18749_ (.A1_N(_09494_),
    .A2_N(_09508_),
    .B1(_09495_),
    .B2(_09489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09637_));
 sky130_fd_sc_hd__a21boi_2 _18750_ (.A1(_09494_),
    .A2(_09508_),
    .B1_N(_09496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09638_));
 sky130_fd_sc_hd__nand2_2 _18751_ (.A(\b_l[5] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09639_));
 sky130_fd_sc_hd__nand2_2 _18752_ (.A(\b_l[3] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09640_));
 sky130_fd_sc_hd__nand2_2 _18753_ (.A(\b_l[4] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09641_));
 sky130_fd_sc_hd__a22oi_2 _18754_ (.A1(\b_l[4] ),
    .A2(\a_l[9] ),
    .B1(\a_l[10] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09642_));
 sky130_fd_sc_hd__nand2_2 _18755_ (.A(_09640_),
    .B(_09641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09643_));
 sky130_fd_sc_hd__and4_2 _18756_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[9] ),
    .D(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09644_));
 sky130_fd_sc_hd__nand4_2 _18757_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[9] ),
    .D(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_2 _18758_ (.A1(_09643_),
    .A2(_09645_),
    .B1(_09639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09647_));
 sky130_fd_sc_hd__o311a_2 _18759_ (.A1(_09275_),
    .A2(_09286_),
    .A3(_04182_),
    .B1(_09639_),
    .C1(_09643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09648_));
 sky130_fd_sc_hd__a41o_2 _18760_ (.A1(\b_l[3] ),
    .A2(\b_l[4] ),
    .A3(\a_l[9] ),
    .A4(\a_l[10] ),
    .B1(_09639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09649_));
 sky130_fd_sc_hd__a22o_2 _18761_ (.A1(\b_l[5] ),
    .A2(\a_l[8] ),
    .B1(_09643_),
    .B2(_09645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09650_));
 sky130_fd_sc_hd__o21ai_2 _18762_ (.A1(_09642_),
    .A2(_09649_),
    .B1(_09650_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09651_));
 sky130_fd_sc_hd__a21oi_2 _18763_ (.A1(_09478_),
    .A2(_09479_),
    .B1(_09487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_2 _18764_ (.A(_09484_),
    .B(_09487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09653_));
 sky130_fd_sc_hd__nand2_2 _18765_ (.A(_09480_),
    .B(_09653_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09654_));
 sky130_fd_sc_hd__nor2_2 _18766_ (.A(_09155_),
    .B(_09297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_2 _18767_ (.A(\b_l[2] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_2 _18768_ (.A(\b_l[0] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09658_));
 sky130_fd_sc_hd__a22oi_2 _18769_ (.A1(\b_l[1] ),
    .A2(\a_l[12] ),
    .B1(\a_l[13] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09659_));
 sky130_fd_sc_hd__nand2_2 _18770_ (.A(_09481_),
    .B(_09658_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09660_));
 sky130_fd_sc_hd__nand4_2 _18771_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[12] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09661_));
 sky130_fd_sc_hd__nand2_2 _18772_ (.A(_09660_),
    .B(_09661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09662_));
 sky130_fd_sc_hd__nand2_2 _18773_ (.A(_09662_),
    .B(_09655_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09663_));
 sky130_fd_sc_hd__o211ai_2 _18774_ (.A1(_09155_),
    .A2(_09297_),
    .B1(_09660_),
    .C1(_09661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09664_));
 sky130_fd_sc_hd__nand4_2 _18775_ (.A(_09660_),
    .B(_09661_),
    .C(\b_l[2] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09665_));
 sky130_fd_sc_hd__o2bb2ai_2 _18776_ (.A1_N(_09660_),
    .A2_N(_09661_),
    .B1(_09155_),
    .B2(_09297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09666_));
 sky130_fd_sc_hd__o211ai_2 _18777_ (.A1(_09483_),
    .A2(_09652_),
    .B1(_09665_),
    .C1(_09666_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09667_));
 sky130_fd_sc_hd__nand3_2 _18778_ (.A(_09663_),
    .B(_09664_),
    .C(_09654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_2 _18779_ (.A(_09667_),
    .B(_09669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09670_));
 sky130_fd_sc_hd__o21ai_2 _18780_ (.A1(_09647_),
    .A2(_09648_),
    .B1(_09670_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09671_));
 sky130_fd_sc_hd__nand3_2 _18781_ (.A(_09651_),
    .B(_09667_),
    .C(_09669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09672_));
 sky130_fd_sc_hd__o211ai_2 _18782_ (.A1(_09647_),
    .A2(_09648_),
    .B1(_09667_),
    .C1(_09669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09673_));
 sky130_fd_sc_hd__nand2_2 _18783_ (.A(_09670_),
    .B(_09651_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09674_));
 sky130_fd_sc_hd__nand2_2 _18784_ (.A(_09671_),
    .B(_09672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09675_));
 sky130_fd_sc_hd__nand3_2 _18785_ (.A(_09674_),
    .B(_09637_),
    .C(_09673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09676_));
 sky130_fd_sc_hd__nand3_2 _18786_ (.A(_09638_),
    .B(_09671_),
    .C(_09672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_2 _18787_ (.A1(_09498_),
    .A2(_09500_),
    .B1(_09502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09678_));
 sky130_fd_sc_hd__nand2_2 _18788_ (.A(\a_l[5] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_2 _18789_ (.A(\a_l[6] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09681_));
 sky130_fd_sc_hd__nand2_2 _18790_ (.A(\b_l[6] ),
    .B(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09682_));
 sky130_fd_sc_hd__a22oi_2 _18791_ (.A1(\b_l[6] ),
    .A2(\a_l[7] ),
    .B1(\b_l[7] ),
    .B2(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09683_));
 sky130_fd_sc_hd__nand2_2 _18792_ (.A(_09681_),
    .B(_09682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09684_));
 sky130_fd_sc_hd__nand4_2 _18793_ (.A(\a_l[6] ),
    .B(\b_l[6] ),
    .C(\a_l[7] ),
    .D(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09685_));
 sky130_fd_sc_hd__nand4_2 _18794_ (.A(_09684_),
    .B(_09685_),
    .C(\a_l[5] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09686_));
 sky130_fd_sc_hd__a22o_2 _18795_ (.A1(\a_l[5] ),
    .A2(\b_l[8] ),
    .B1(_09684_),
    .B2(_09685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09687_));
 sky130_fd_sc_hd__nand3_2 _18796_ (.A(_09687_),
    .B(_09678_),
    .C(_09686_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09688_));
 sky130_fd_sc_hd__o211ai_2 _18797_ (.A1(_09210_),
    .A2(_09264_),
    .B1(_09684_),
    .C1(_09685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09689_));
 sky130_fd_sc_hd__a21o_2 _18798_ (.A1(_09684_),
    .A2(_09685_),
    .B1(_09680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09691_));
 sky130_fd_sc_hd__nand3b_2 _18799_ (.A_N(_09678_),
    .B(_09689_),
    .C(_09691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09692_));
 sky130_fd_sc_hd__nand2_2 _18800_ (.A(_09688_),
    .B(_09692_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09693_));
 sky130_fd_sc_hd__a32o_2 _18801_ (.A1(\a_l[5] ),
    .A2(\a_l[6] ),
    .A3(_04259_),
    .B1(_09454_),
    .B2(_09451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09694_));
 sky130_fd_sc_hd__and2_2 _18802_ (.A(_09693_),
    .B(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09695_));
 sky130_fd_sc_hd__nor2_2 _18803_ (.A(_09694_),
    .B(_09693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09696_));
 sky130_fd_sc_hd__a21oi_2 _18804_ (.A1(_09688_),
    .A2(_09692_),
    .B1(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09697_));
 sky130_fd_sc_hd__a21o_2 _18805_ (.A1(_09688_),
    .A2(_09692_),
    .B1(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09698_));
 sky130_fd_sc_hd__nand2_2 _18806_ (.A(_09692_),
    .B(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09699_));
 sky130_fd_sc_hd__and3_2 _18807_ (.A(_09688_),
    .B(_09692_),
    .C(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09700_));
 sky130_fd_sc_hd__nand3_2 _18808_ (.A(_09688_),
    .B(_09692_),
    .C(_09694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09701_));
 sky130_fd_sc_hd__o2bb2ai_2 _18809_ (.A1_N(_09676_),
    .A2_N(_09677_),
    .B1(_09695_),
    .B2(_09696_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09702_));
 sky130_fd_sc_hd__o21ai_2 _18810_ (.A1(_09697_),
    .A2(_09700_),
    .B1(_09676_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09703_));
 sky130_fd_sc_hd__o211ai_2 _18811_ (.A1(_09697_),
    .A2(_09700_),
    .B1(_09676_),
    .C1(_09677_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09704_));
 sky130_fd_sc_hd__nand4_2 _18812_ (.A(_09676_),
    .B(_09677_),
    .C(_09698_),
    .D(_09701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09705_));
 sky130_fd_sc_hd__o2bb2ai_2 _18813_ (.A1_N(_09676_),
    .A2_N(_09677_),
    .B1(_09697_),
    .B2(_09700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09706_));
 sky130_fd_sc_hd__o211ai_2 _18814_ (.A1(_09511_),
    .A2(_09520_),
    .B1(_09705_),
    .C1(_09706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09707_));
 sky130_fd_sc_hd__nand3_2 _18815_ (.A(_09702_),
    .B(_09704_),
    .C(_09636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09708_));
 sky130_fd_sc_hd__nand2_2 _18816_ (.A(_09707_),
    .B(_09708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09709_));
 sky130_fd_sc_hd__nand4_2 _18817_ (.A(_09632_),
    .B(_09633_),
    .C(_09707_),
    .D(_09708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09710_));
 sky130_fd_sc_hd__nand2_2 _18818_ (.A(_09709_),
    .B(_09634_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09711_));
 sky130_fd_sc_hd__nand4_2 _18819_ (.A(_09630_),
    .B(_09631_),
    .C(_09707_),
    .D(_09708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09712_));
 sky130_fd_sc_hd__a22o_2 _18820_ (.A1(_09630_),
    .A2(_09631_),
    .B1(_09707_),
    .B2(_09708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09713_));
 sky130_fd_sc_hd__a21oi_2 _18821_ (.A1(_09530_),
    .A2(_09562_),
    .B1(_09528_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09714_));
 sky130_fd_sc_hd__o2bb2ai_2 _18822_ (.A1_N(_09562_),
    .A2_N(_09530_),
    .B1(_09527_),
    .B2(_09522_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09715_));
 sky130_fd_sc_hd__nand3_2 _18823_ (.A(_09712_),
    .B(_09713_),
    .C(_09715_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09716_));
 sky130_fd_sc_hd__nand3_2 _18824_ (.A(_09714_),
    .B(_09711_),
    .C(_09710_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09717_));
 sky130_fd_sc_hd__a31o_2 _18825_ (.A1(_09547_),
    .A2(_09550_),
    .A3(_09551_),
    .B1(_09556_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09718_));
 sky130_fd_sc_hd__a21oi_2 _18826_ (.A1(_09716_),
    .A2(_09717_),
    .B1(_09718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09719_));
 sky130_fd_sc_hd__a21o_2 _18827_ (.A1(_09716_),
    .A2(_09717_),
    .B1(_09718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09720_));
 sky130_fd_sc_hd__o211a_2 _18828_ (.A1(_09554_),
    .A2(_09556_),
    .B1(_09716_),
    .C1(_09717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09721_));
 sky130_fd_sc_hd__o211ai_2 _18829_ (.A1(_09554_),
    .A2(_09556_),
    .B1(_09716_),
    .C1(_09717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09722_));
 sky130_fd_sc_hd__nand2_2 _18830_ (.A(_09572_),
    .B(_09416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09723_));
 sky130_fd_sc_hd__o2bb2ai_2 _18831_ (.A1_N(_09416_),
    .A2_N(_09572_),
    .B1(_09573_),
    .B2(_09565_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09724_));
 sky130_fd_sc_hd__o21bai_2 _18832_ (.A1(_09719_),
    .A2(_09721_),
    .B1_N(_09724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09725_));
 sky130_fd_sc_hd__a21oi_2 _18833_ (.A1(_09574_),
    .A2(_09723_),
    .B1(_09719_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09726_));
 sky130_fd_sc_hd__nand3_2 _18834_ (.A(_09720_),
    .B(_09722_),
    .C(_09724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09727_));
 sky130_fd_sc_hd__a21oi_2 _18835_ (.A1(_09725_),
    .A2(_09727_),
    .B1(_09582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09728_));
 sky130_fd_sc_hd__a21oi_2 _18836_ (.A1(_09726_),
    .A2(_09722_),
    .B1(_09583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09729_));
 sky130_fd_sc_hd__nand2_2 _18837_ (.A(_09729_),
    .B(_09725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09730_));
 sky130_fd_sc_hd__a21oi_2 _18838_ (.A1(_09725_),
    .A2(_09729_),
    .B1(_09728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09731_));
 sky130_fd_sc_hd__a2bb2o_2 _18839_ (.A1_N(_09588_),
    .A2_N(_09591_),
    .B1(_09580_),
    .B2(_09586_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09732_));
 sky130_fd_sc_hd__or3_2 _18840_ (.A(_09437_),
    .B(_09584_),
    .C(_09728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09733_));
 sky130_fd_sc_hd__o2111ai_2 _18841_ (.A1(_09313_),
    .A2(_09438_),
    .B1(_09587_),
    .C1(_09731_),
    .D1(_09590_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09734_));
 sky130_fd_sc_hd__o31a_2 _18842_ (.A1(_09437_),
    .A2(_09584_),
    .A3(_09728_),
    .B1(_09734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09735_));
 sky130_fd_sc_hd__o211a_2 _18843_ (.A1(_09731_),
    .A2(_09732_),
    .B1(_09735_),
    .C1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00383_));
 sky130_fd_sc_hd__o211a_2 _18844_ (.A1(_09625_),
    .A2(_09629_),
    .B1(_05043_),
    .C1(_06401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09736_));
 sky130_fd_sc_hd__a211o_2 _18845_ (.A1(_09626_),
    .A2(_09630_),
    .B1(_05044_),
    .C1(_06402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09737_));
 sky130_fd_sc_hd__o311a_2 _18846_ (.A1(_09329_),
    .A2(_09351_),
    .A3(_06402_),
    .B1(_09626_),
    .C1(_09630_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09738_));
 sky130_fd_sc_hd__nor2_2 _18847_ (.A(_09736_),
    .B(_09738_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09739_));
 sky130_fd_sc_hd__a21boi_2 _18848_ (.A1(_09619_),
    .A2(_09598_),
    .B1_N(_09612_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09740_));
 sky130_fd_sc_hd__nand2_2 _18849_ (.A(_09688_),
    .B(_09699_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09741_));
 sky130_fd_sc_hd__a21boi_2 _18850_ (.A1(_09692_),
    .A2(_09694_),
    .B1_N(_09688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09742_));
 sky130_fd_sc_hd__a22o_2 _18851_ (.A1(\a_l[2] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09743_));
 sky130_fd_sc_hd__nand4_2 _18852_ (.A(\a_l[2] ),
    .B(\a_l[1] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09744_));
 sky130_fd_sc_hd__o2111ai_2 _18853_ (.A1(_05044_),
    .A2(_06441_),
    .B1(\a_l[0] ),
    .C1(\b_l[14] ),
    .D1(_09743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09745_));
 sky130_fd_sc_hd__a22o_2 _18854_ (.A1(\a_l[0] ),
    .A2(\b_l[14] ),
    .B1(_09743_),
    .B2(_09744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09746_));
 sky130_fd_sc_hd__nand2_2 _18855_ (.A(_09745_),
    .B(_09746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09747_));
 sky130_fd_sc_hd__a21oi_2 _18856_ (.A1(_09603_),
    .A2(_09604_),
    .B1(_09609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_2 _18857_ (.A(\a_l[3] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_2 _18858_ (.A(\a_l[4] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09750_));
 sky130_fd_sc_hd__nand2_2 _18859_ (.A(\a_l[5] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09751_));
 sky130_fd_sc_hd__a22oi_2 _18860_ (.A1(\a_l[5] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_2 _18861_ (.A(_09750_),
    .B(_09751_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09753_));
 sky130_fd_sc_hd__nand4_2 _18862_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09754_));
 sky130_fd_sc_hd__a22oi_2 _18863_ (.A1(\a_l[3] ),
    .A2(\b_l[11] ),
    .B1(_09753_),
    .B2(_09754_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09755_));
 sky130_fd_sc_hd__a21bo_2 _18864_ (.A1(_09753_),
    .A2(_09754_),
    .B1_N(_09749_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09756_));
 sky130_fd_sc_hd__o2111a_2 _18865_ (.A1(_04555_),
    .A2(_06605_),
    .B1(\a_l[3] ),
    .C1(\b_l[11] ),
    .D1(_09753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09757_));
 sky130_fd_sc_hd__o2111ai_2 _18866_ (.A1(_04555_),
    .A2(_06605_),
    .B1(\a_l[3] ),
    .C1(\b_l[11] ),
    .D1(_09753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09758_));
 sky130_fd_sc_hd__o22a_2 _18867_ (.A1(_09605_),
    .A2(_09616_),
    .B1(_09755_),
    .B2(_09757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09759_));
 sky130_fd_sc_hd__o22ai_2 _18868_ (.A1(_09605_),
    .A2(_09616_),
    .B1(_09755_),
    .B2(_09757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09760_));
 sky130_fd_sc_hd__o211ai_2 _18869_ (.A1(_09607_),
    .A2(_09748_),
    .B1(_09756_),
    .C1(_09758_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09761_));
 sky130_fd_sc_hd__a21o_2 _18870_ (.A1(_09760_),
    .A2(_09761_),
    .B1(_09747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09762_));
 sky130_fd_sc_hd__nand3_2 _18871_ (.A(_09747_),
    .B(_09760_),
    .C(_09761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09763_));
 sky130_fd_sc_hd__nand4_2 _18872_ (.A(_09745_),
    .B(_09746_),
    .C(_09760_),
    .D(_09761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09764_));
 sky130_fd_sc_hd__a22o_2 _18873_ (.A1(_09745_),
    .A2(_09746_),
    .B1(_09760_),
    .B2(_09761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09765_));
 sky130_fd_sc_hd__nand3_2 _18874_ (.A(_09765_),
    .B(_09741_),
    .C(_09764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09766_));
 sky130_fd_sc_hd__nand3_2 _18875_ (.A(_09742_),
    .B(_09762_),
    .C(_09763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09767_));
 sky130_fd_sc_hd__a31o_2 _18876_ (.A1(_09742_),
    .A2(_09762_),
    .A3(_09763_),
    .B1(_09740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09768_));
 sky130_fd_sc_hd__a22o_2 _18877_ (.A1(_09612_),
    .A2(_09621_),
    .B1(_09766_),
    .B2(_09767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09769_));
 sky130_fd_sc_hd__nand4_2 _18878_ (.A(_09612_),
    .B(_09621_),
    .C(_09766_),
    .D(_09767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09770_));
 sky130_fd_sc_hd__nand2_2 _18879_ (.A(_09769_),
    .B(_09770_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09771_));
 sky130_fd_sc_hd__nand2_2 _18880_ (.A(_09677_),
    .B(_09703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09772_));
 sky130_fd_sc_hd__o21a_2 _18881_ (.A1(_09637_),
    .A2(_09675_),
    .B1(_09703_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09773_));
 sky130_fd_sc_hd__a21oi_2 _18882_ (.A1(_09640_),
    .A2(_09641_),
    .B1(_09639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09774_));
 sky130_fd_sc_hd__a21o_2 _18883_ (.A1(_09639_),
    .A2(_09645_),
    .B1(_09642_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09775_));
 sky130_fd_sc_hd__nand2_2 _18884_ (.A(\a_l[6] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_2 _18885_ (.A(\a_l[7] ),
    .B(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_2 _18886_ (.A(\b_l[6] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09778_));
 sky130_fd_sc_hd__nand2_2 _18887_ (.A(_09777_),
    .B(_09778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09779_));
 sky130_fd_sc_hd__nand4_2 _18888_ (.A(\b_l[6] ),
    .B(\a_l[7] ),
    .C(\b_l[7] ),
    .D(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09780_));
 sky130_fd_sc_hd__a21o_2 _18889_ (.A1(_09779_),
    .A2(_09780_),
    .B1(_09776_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09781_));
 sky130_fd_sc_hd__o211ai_2 _18890_ (.A1(_09231_),
    .A2(_09264_),
    .B1(_09779_),
    .C1(_09780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09782_));
 sky130_fd_sc_hd__nand4_2 _18891_ (.A(_09779_),
    .B(_09780_),
    .C(\a_l[6] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09783_));
 sky130_fd_sc_hd__a22o_2 _18892_ (.A1(\a_l[6] ),
    .A2(\b_l[8] ),
    .B1(_09779_),
    .B2(_09780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09784_));
 sky130_fd_sc_hd__a21oi_2 _18893_ (.A1(_09781_),
    .A2(_09782_),
    .B1(_09775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09785_));
 sky130_fd_sc_hd__o211ai_2 _18894_ (.A1(_09644_),
    .A2(_09774_),
    .B1(_09783_),
    .C1(_09784_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09786_));
 sky130_fd_sc_hd__nand3_2 _18895_ (.A(_09781_),
    .B(_09782_),
    .C(_09775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09787_));
 sky130_fd_sc_hd__o21ai_2 _18896_ (.A1(_09680_),
    .A2(_09683_),
    .B1(_09685_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09788_));
 sky130_fd_sc_hd__a21bo_2 _18897_ (.A1(_09786_),
    .A2(_09787_),
    .B1_N(_09788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09789_));
 sky130_fd_sc_hd__o2111ai_2 _18898_ (.A1(_09680_),
    .A2(_09683_),
    .B1(_09685_),
    .C1(_09786_),
    .D1(_09787_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09790_));
 sky130_fd_sc_hd__a21o_2 _18899_ (.A1(_09786_),
    .A2(_09787_),
    .B1(_09788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09791_));
 sky130_fd_sc_hd__nand3_2 _18900_ (.A(_09786_),
    .B(_09787_),
    .C(_09788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_2 _18901_ (.A(_09791_),
    .B(_09792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_2 _18902_ (.A(_09789_),
    .B(_09790_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_2 _18903_ (.A(_09651_),
    .B(_09667_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_2 _18904_ (.A(_09669_),
    .B(_09795_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09796_));
 sky130_fd_sc_hd__a21boi_2 _18905_ (.A1(_09651_),
    .A2(_09667_),
    .B1_N(_09669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09797_));
 sky130_fd_sc_hd__nand2_2 _18906_ (.A(\b_l[5] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09798_));
 sky130_fd_sc_hd__a22oi_2 _18907_ (.A1(\b_l[4] ),
    .A2(\a_l[10] ),
    .B1(\a_l[11] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09799_));
 sky130_fd_sc_hd__and4_2 _18908_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[10] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09800_));
 sky130_fd_sc_hd__nand4_2 _18909_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[10] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09801_));
 sky130_fd_sc_hd__o21ai_2 _18910_ (.A1(_09799_),
    .A2(_09800_),
    .B1(_09798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09802_));
 sky130_fd_sc_hd__nand4b_2 _18911_ (.A_N(_09799_),
    .B(_09801_),
    .C(\b_l[5] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09803_));
 sky130_fd_sc_hd__o21bai_2 _18912_ (.A1(_09799_),
    .A2(_09800_),
    .B1_N(_09798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09804_));
 sky130_fd_sc_hd__o21a_2 _18913_ (.A1(_09220_),
    .A2(_09275_),
    .B1(_09801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09805_));
 sky130_fd_sc_hd__o21ai_2 _18914_ (.A1(_09220_),
    .A2(_09275_),
    .B1(_09801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09806_));
 sky130_fd_sc_hd__o21ai_2 _18915_ (.A1(_09799_),
    .A2(_09806_),
    .B1(_09804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09807_));
 sky130_fd_sc_hd__nand2_2 _18916_ (.A(_09802_),
    .B(_09803_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09808_));
 sky130_fd_sc_hd__a21o_2 _18917_ (.A1(_09656_),
    .A2(_09661_),
    .B1(_09659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09809_));
 sky130_fd_sc_hd__a21oi_2 _18918_ (.A1(_09656_),
    .A2(_09661_),
    .B1(_09659_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09810_));
 sky130_fd_sc_hd__nand2_2 _18919_ (.A(\b_l[2] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_2 _18920_ (.A(\b_l[1] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_2 _18921_ (.A(\b_l[0] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09813_));
 sky130_fd_sc_hd__a22oi_2 _18922_ (.A1(\b_l[1] ),
    .A2(\a_l[13] ),
    .B1(\a_l[14] ),
    .B2(\b_l[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_2 _18923_ (.A(_09812_),
    .B(_09813_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_2 _18924_ (.A(\b_l[1] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09816_));
 sky130_fd_sc_hd__nand4_2 _18925_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[13] ),
    .D(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09817_));
 sky130_fd_sc_hd__o2bb2ai_2 _18926_ (.A1_N(_09815_),
    .A2_N(_09817_),
    .B1(_09155_),
    .B2(_09319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09818_));
 sky130_fd_sc_hd__nand3_2 _18927_ (.A(_09817_),
    .B(\a_l[12] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09819_));
 sky130_fd_sc_hd__o221a_2 _18928_ (.A1(_09155_),
    .A2(_09319_),
    .B1(_09658_),
    .B2(_09816_),
    .C1(_09815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09820_));
 sky130_fd_sc_hd__o221ai_2 _18929_ (.A1(_09155_),
    .A2(_09319_),
    .B1(_09658_),
    .B2(_09816_),
    .C1(_09815_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09821_));
 sky130_fd_sc_hd__a21o_2 _18930_ (.A1(_09815_),
    .A2(_09817_),
    .B1(_09811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09822_));
 sky130_fd_sc_hd__nand2_2 _18931_ (.A(_09822_),
    .B(_09809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09823_));
 sky130_fd_sc_hd__nand3_2 _18932_ (.A(_09822_),
    .B(_09809_),
    .C(_09821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09824_));
 sky130_fd_sc_hd__o211a_2 _18933_ (.A1(_09819_),
    .A2(_09814_),
    .B1(_09810_),
    .C1(_09818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09825_));
 sky130_fd_sc_hd__o211ai_2 _18934_ (.A1(_09819_),
    .A2(_09814_),
    .B1(_09810_),
    .C1(_09818_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_2 _18935_ (.A(_09824_),
    .B(_09826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09827_));
 sky130_fd_sc_hd__and3_2 _18936_ (.A(_09808_),
    .B(_09824_),
    .C(_09826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09828_));
 sky130_fd_sc_hd__o2111ai_2 _18937_ (.A1(_09806_),
    .A2(_09799_),
    .B1(_09804_),
    .C1(_09824_),
    .D1(_09826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09829_));
 sky130_fd_sc_hd__nand2_2 _18938_ (.A(_09827_),
    .B(_09807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09830_));
 sky130_fd_sc_hd__nand2_2 _18939_ (.A(_09807_),
    .B(_09824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09831_));
 sky130_fd_sc_hd__and3_2 _18940_ (.A(_09826_),
    .B(_09807_),
    .C(_09824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09832_));
 sky130_fd_sc_hd__a21o_2 _18941_ (.A1(_09824_),
    .A2(_09826_),
    .B1(_09807_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09833_));
 sky130_fd_sc_hd__nand2_2 _18942_ (.A(_09796_),
    .B(_09830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09834_));
 sky130_fd_sc_hd__nand3_2 _18943_ (.A(_09796_),
    .B(_09829_),
    .C(_09830_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09835_));
 sky130_fd_sc_hd__nand2_2 _18944_ (.A(_09797_),
    .B(_09833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09836_));
 sky130_fd_sc_hd__o211ai_2 _18945_ (.A1(_09831_),
    .A2(_09825_),
    .B1(_09797_),
    .C1(_09833_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09837_));
 sky130_fd_sc_hd__o221ai_2 _18946_ (.A1(_09828_),
    .A2(_09834_),
    .B1(_09832_),
    .B2(_09836_),
    .C1(_09793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09838_));
 sky130_fd_sc_hd__a22o_2 _18947_ (.A1(_09789_),
    .A2(_09790_),
    .B1(_09835_),
    .B2(_09837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09839_));
 sky130_fd_sc_hd__and3_2 _18948_ (.A(_09794_),
    .B(_09835_),
    .C(_09837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09840_));
 sky130_fd_sc_hd__nand4_2 _18949_ (.A(_09791_),
    .B(_09792_),
    .C(_09835_),
    .D(_09837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09841_));
 sky130_fd_sc_hd__a22o_2 _18950_ (.A1(_09791_),
    .A2(_09792_),
    .B1(_09835_),
    .B2(_09837_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09842_));
 sky130_fd_sc_hd__nand2_2 _18951_ (.A(_09773_),
    .B(_09842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09843_));
 sky130_fd_sc_hd__nand3_2 _18952_ (.A(_09773_),
    .B(_09841_),
    .C(_09842_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09844_));
 sky130_fd_sc_hd__nand3_2 _18953_ (.A(_09839_),
    .B(_09772_),
    .C(_09838_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09845_));
 sky130_fd_sc_hd__a22o_2 _18954_ (.A1(_09769_),
    .A2(_09770_),
    .B1(_09844_),
    .B2(_09845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09846_));
 sky130_fd_sc_hd__nand4_2 _18955_ (.A(_09769_),
    .B(_09770_),
    .C(_09844_),
    .D(_09845_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09847_));
 sky130_fd_sc_hd__a21o_2 _18956_ (.A1(_09844_),
    .A2(_09845_),
    .B1(_09771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09848_));
 sky130_fd_sc_hd__o211ai_2 _18957_ (.A1(_09840_),
    .A2(_09843_),
    .B1(_09845_),
    .C1(_09771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09849_));
 sky130_fd_sc_hd__nand2_2 _18958_ (.A(_09848_),
    .B(_09849_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09850_));
 sky130_fd_sc_hd__a21boi_2 _18959_ (.A1(_09634_),
    .A2(_09708_),
    .B1_N(_09707_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09851_));
 sky130_fd_sc_hd__nand3_2 _18960_ (.A(_09846_),
    .B(_09847_),
    .C(_09851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09852_));
 sky130_fd_sc_hd__nand3b_2 _18961_ (.A_N(_09851_),
    .B(_09849_),
    .C(_09848_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09853_));
 sky130_fd_sc_hd__o221ai_2 _18962_ (.A1(_09736_),
    .A2(_09738_),
    .B1(_09851_),
    .B2(_09850_),
    .C1(_09852_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09854_));
 sky130_fd_sc_hd__a21bo_2 _18963_ (.A1(_09852_),
    .A2(_09853_),
    .B1_N(_09739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09855_));
 sky130_fd_sc_hd__nand4_2 _18964_ (.A(_09716_),
    .B(_09722_),
    .C(_09854_),
    .D(_09855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09856_));
 sky130_fd_sc_hd__a22oi_2 _18965_ (.A1(_09716_),
    .A2(_09722_),
    .B1(_09854_),
    .B2(_09855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09857_));
 sky130_fd_sc_hd__a22o_2 _18966_ (.A1(_09716_),
    .A2(_09722_),
    .B1(_09854_),
    .B2(_09855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09858_));
 sky130_fd_sc_hd__nand2_2 _18967_ (.A(_09856_),
    .B(_09858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09859_));
 sky130_fd_sc_hd__a22oi_2 _18968_ (.A1(_09726_),
    .A2(_09722_),
    .B1(_09858_),
    .B2(_09856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09860_));
 sky130_fd_sc_hd__and4_2 _18969_ (.A(_09722_),
    .B(_09858_),
    .C(_09726_),
    .D(_09856_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09861_));
 sky130_fd_sc_hd__or2_2 _18970_ (.A(_09860_),
    .B(_09861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09862_));
 sky130_fd_sc_hd__a21oi_2 _18971_ (.A1(_09730_),
    .A2(_09735_),
    .B1(_09862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09863_));
 sky130_fd_sc_hd__a31o_2 _18972_ (.A1(_09730_),
    .A2(_09735_),
    .A3(_09862_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09864_));
 sky130_fd_sc_hd__nor2_2 _18973_ (.A(_09863_),
    .B(_09864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00384_));
 sky130_fd_sc_hd__nor2_2 _18974_ (.A(_09861_),
    .B(_09863_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_2 _18975_ (.A(_09852_),
    .B(_09739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09866_));
 sky130_fd_sc_hd__o21ai_2 _18976_ (.A1(_09850_),
    .A2(_09851_),
    .B1(_09866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09867_));
 sky130_fd_sc_hd__a21boi_2 _18977_ (.A1(_09739_),
    .A2(_09852_),
    .B1_N(_09853_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09868_));
 sky130_fd_sc_hd__o2bb2ai_2 _18978_ (.A1_N(_09771_),
    .A2_N(_09845_),
    .B1(_09843_),
    .B2(_09840_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09869_));
 sky130_fd_sc_hd__a21boi_2 _18979_ (.A1(_09771_),
    .A2(_09845_),
    .B1_N(_09844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09870_));
 sky130_fd_sc_hd__a21o_2 _18980_ (.A1(_09787_),
    .A2(_09788_),
    .B1(_09785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09871_));
 sky130_fd_sc_hd__a21oi_2 _18981_ (.A1(_09787_),
    .A2(_09788_),
    .B1(_09785_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09872_));
 sky130_fd_sc_hd__a22o_2 _18982_ (.A1(\a_l[3] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09873_));
 sky130_fd_sc_hd__and3_2 _18983_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09874_));
 sky130_fd_sc_hd__nand4_2 _18984_ (.A(\a_l[2] ),
    .B(\a_l[3] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09875_));
 sky130_fd_sc_hd__and3_2 _18985_ (.A(_09875_),
    .B(\b_l[14] ),
    .C(\a_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09876_));
 sky130_fd_sc_hd__and4_2 _18986_ (.A(_09873_),
    .B(_09875_),
    .C(\a_l[1] ),
    .D(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09877_));
 sky130_fd_sc_hd__a22oi_2 _18987_ (.A1(\a_l[1] ),
    .A2(\b_l[14] ),
    .B1(_09873_),
    .B2(_09875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09878_));
 sky130_fd_sc_hd__a21oi_2 _18988_ (.A1(_09873_),
    .A2(_09876_),
    .B1(_09878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09879_));
 sky130_fd_sc_hd__a21o_2 _18989_ (.A1(_09749_),
    .A2(_09754_),
    .B1(_09752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09880_));
 sky130_fd_sc_hd__a21oi_2 _18990_ (.A1(_09749_),
    .A2(_09754_),
    .B1(_09752_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09881_));
 sky130_fd_sc_hd__nand2_2 _18991_ (.A(\a_l[5] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09882_));
 sky130_fd_sc_hd__nand2_2 _18992_ (.A(\a_l[6] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09883_));
 sky130_fd_sc_hd__a22oi_2 _18993_ (.A1(\a_l[6] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09884_));
 sky130_fd_sc_hd__nand2_2 _18994_ (.A(_09882_),
    .B(_09883_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09885_));
 sky130_fd_sc_hd__nand4_2 _18995_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09886_));
 sky130_fd_sc_hd__nand2_2 _18996_ (.A(\a_l[4] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09887_));
 sky130_fd_sc_hd__a21o_2 _18997_ (.A1(_09885_),
    .A2(_09886_),
    .B1(_09887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09888_));
 sky130_fd_sc_hd__o21ai_2 _18998_ (.A1(_09882_),
    .A2(_09883_),
    .B1(_09887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09889_));
 sky130_fd_sc_hd__o211ai_2 _18999_ (.A1(_09884_),
    .A2(_09889_),
    .B1(_09880_),
    .C1(_09888_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09890_));
 sky130_fd_sc_hd__nand3_2 _19000_ (.A(_09886_),
    .B(\b_l[11] ),
    .C(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09891_));
 sky130_fd_sc_hd__o2bb2ai_2 _19001_ (.A1_N(_09885_),
    .A2_N(_09886_),
    .B1(_09199_),
    .B2(_09308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09892_));
 sky130_fd_sc_hd__o211a_2 _19002_ (.A1(_09891_),
    .A2(_09884_),
    .B1(_09881_),
    .C1(_09892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09893_));
 sky130_fd_sc_hd__o211ai_2 _19003_ (.A1(_09891_),
    .A2(_09884_),
    .B1(_09881_),
    .C1(_09892_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09894_));
 sky130_fd_sc_hd__nand2_2 _19004_ (.A(_09890_),
    .B(_09894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09895_));
 sky130_fd_sc_hd__o21ai_2 _19005_ (.A1(_09877_),
    .A2(_09878_),
    .B1(_09895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09896_));
 sky130_fd_sc_hd__nand2_2 _19006_ (.A(_09879_),
    .B(_09890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09897_));
 sky130_fd_sc_hd__o211ai_2 _19007_ (.A1(_09877_),
    .A2(_09878_),
    .B1(_09890_),
    .C1(_09894_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09898_));
 sky130_fd_sc_hd__nand2_2 _19008_ (.A(_09895_),
    .B(_09879_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09899_));
 sky130_fd_sc_hd__nand3_2 _19009_ (.A(_09872_),
    .B(_09898_),
    .C(_09899_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09900_));
 sky130_fd_sc_hd__o211ai_2 _19010_ (.A1(_09893_),
    .A2(_09897_),
    .B1(_09896_),
    .C1(_09871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09901_));
 sky130_fd_sc_hd__o41a_2 _19011_ (.A1(_09605_),
    .A2(_09616_),
    .A3(_09755_),
    .A4(_09757_),
    .B1(_09747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09902_));
 sky130_fd_sc_hd__nand2_2 _19012_ (.A(_09747_),
    .B(_09761_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09903_));
 sky130_fd_sc_hd__nand4_2 _19013_ (.A(_09760_),
    .B(_09900_),
    .C(_09901_),
    .D(_09903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09904_));
 sky130_fd_sc_hd__o2bb2ai_2 _19014_ (.A1_N(_09900_),
    .A2_N(_09901_),
    .B1(_09902_),
    .B2(_09759_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09905_));
 sky130_fd_sc_hd__nand2_2 _19015_ (.A(_09904_),
    .B(_09905_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09906_));
 sky130_fd_sc_hd__and2_2 _19016_ (.A(\a_l[7] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09907_));
 sky130_fd_sc_hd__nand2_2 _19017_ (.A(\b_l[7] ),
    .B(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_2 _19018_ (.A(\b_l[6] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09909_));
 sky130_fd_sc_hd__nand2_2 _19019_ (.A(_09908_),
    .B(_09909_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09910_));
 sky130_fd_sc_hd__nand4_2 _19020_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[8] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09911_));
 sky130_fd_sc_hd__a21oi_2 _19021_ (.A1(_09910_),
    .A2(_09911_),
    .B1(_09907_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09912_));
 sky130_fd_sc_hd__a22o_2 _19022_ (.A1(\a_l[7] ),
    .A2(\b_l[8] ),
    .B1(_09910_),
    .B2(_09911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09913_));
 sky130_fd_sc_hd__o211a_2 _19023_ (.A1(_04260_),
    .A2(_06985_),
    .B1(_09907_),
    .C1(_09910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09914_));
 sky130_fd_sc_hd__o2111ai_2 _19024_ (.A1(_04260_),
    .A2(_06985_),
    .B1(\a_l[7] ),
    .C1(\b_l[8] ),
    .D1(_09910_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09915_));
 sky130_fd_sc_hd__o21ai_2 _19025_ (.A1(_09798_),
    .A2(_09799_),
    .B1(_09801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09916_));
 sky130_fd_sc_hd__o22ai_2 _19026_ (.A1(_09799_),
    .A2(_09805_),
    .B1(_09912_),
    .B2(_09914_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09917_));
 sky130_fd_sc_hd__nand3_2 _19027_ (.A(_09913_),
    .B(_09915_),
    .C(_09916_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09918_));
 sky130_fd_sc_hd__nand2_2 _19028_ (.A(_09917_),
    .B(_09918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09919_));
 sky130_fd_sc_hd__a21boi_2 _19029_ (.A1(_09776_),
    .A2(_09780_),
    .B1_N(_09779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_2 _19030_ (.A(_09917_),
    .B(_09920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09921_));
 sky130_fd_sc_hd__nand2_2 _19031_ (.A(_09919_),
    .B(_09920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09922_));
 sky130_fd_sc_hd__nand3b_2 _19032_ (.A_N(_09920_),
    .B(_09918_),
    .C(_09917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_2 _19033_ (.A(_09922_),
    .B(_09923_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09924_));
 sky130_fd_sc_hd__o2bb2ai_2 _19034_ (.A1_N(_09808_),
    .A2_N(_09826_),
    .B1(_09823_),
    .B2(_09820_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_2 _19035_ (.A(_09826_),
    .B(_09831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09926_));
 sky130_fd_sc_hd__a21o_2 _19036_ (.A1(_09811_),
    .A2(_09817_),
    .B1(_09814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09927_));
 sky130_fd_sc_hd__a21oi_2 _19037_ (.A1(_09811_),
    .A2(_09817_),
    .B1(_09814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_2 _19038_ (.A(\b_l[2] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09929_));
 sky130_fd_sc_hd__nand2_2 _19039_ (.A(\b_l[0] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_2 _19040_ (.A(_09816_),
    .B(_09930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09931_));
 sky130_fd_sc_hd__nand4_2 _19041_ (.A(\b_l[0] ),
    .B(\b_l[1] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09932_));
 sky130_fd_sc_hd__o211ai_2 _19042_ (.A1(_09155_),
    .A2(_09340_),
    .B1(_09931_),
    .C1(_09932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09933_));
 sky130_fd_sc_hd__a21o_2 _19043_ (.A1(_09931_),
    .A2(_09932_),
    .B1(_09929_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09934_));
 sky130_fd_sc_hd__o2bb2ai_2 _19044_ (.A1_N(_09931_),
    .A2_N(_09932_),
    .B1(_09155_),
    .B2(_09340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09935_));
 sky130_fd_sc_hd__nand4_2 _19045_ (.A(_09931_),
    .B(_09932_),
    .C(\b_l[2] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09936_));
 sky130_fd_sc_hd__nand3_2 _19046_ (.A(_09934_),
    .B(_09927_),
    .C(_09933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09937_));
 sky130_fd_sc_hd__nand3_2 _19047_ (.A(_09928_),
    .B(_09935_),
    .C(_09936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09938_));
 sky130_fd_sc_hd__nand2_2 _19048_ (.A(\b_l[5] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09939_));
 sky130_fd_sc_hd__a22oi_2 _19049_ (.A1(\b_l[4] ),
    .A2(\a_l[11] ),
    .B1(\a_l[12] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09940_));
 sky130_fd_sc_hd__a22o_2 _19050_ (.A1(\b_l[4] ),
    .A2(\a_l[11] ),
    .B1(\a_l[12] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09941_));
 sky130_fd_sc_hd__nand2_2 _19051_ (.A(\b_l[4] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09942_));
 sky130_fd_sc_hd__nand4_2 _19052_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[11] ),
    .D(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09943_));
 sky130_fd_sc_hd__o2bb2a_2 _19053_ (.A1_N(_09941_),
    .A2_N(_09943_),
    .B1(_09220_),
    .B2(_09286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09944_));
 sky130_fd_sc_hd__and4_2 _19054_ (.A(_09941_),
    .B(_09943_),
    .C(\b_l[5] ),
    .D(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09945_));
 sky130_fd_sc_hd__nand2_2 _19055_ (.A(_09939_),
    .B(_09943_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09946_));
 sky130_fd_sc_hd__nor2_2 _19056_ (.A(_09940_),
    .B(_09946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09947_));
 sky130_fd_sc_hd__a21oi_2 _19057_ (.A1(_09941_),
    .A2(_09943_),
    .B1(_09939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09948_));
 sky130_fd_sc_hd__nor2_2 _19058_ (.A(_09947_),
    .B(_09948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09949_));
 sky130_fd_sc_hd__o2bb2ai_2 _19059_ (.A1_N(_09937_),
    .A2_N(_09938_),
    .B1(_09947_),
    .B2(_09948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09950_));
 sky130_fd_sc_hd__nand2_2 _19060_ (.A(_09938_),
    .B(_09949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09951_));
 sky130_fd_sc_hd__nand3_2 _19061_ (.A(_09937_),
    .B(_09938_),
    .C(_09949_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09952_));
 sky130_fd_sc_hd__o211a_2 _19062_ (.A1(_09947_),
    .A2(_09948_),
    .B1(_09937_),
    .C1(_09938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09953_));
 sky130_fd_sc_hd__o211ai_2 _19063_ (.A1(_09947_),
    .A2(_09948_),
    .B1(_09937_),
    .C1(_09938_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09954_));
 sky130_fd_sc_hd__o2bb2ai_2 _19064_ (.A1_N(_09937_),
    .A2_N(_09938_),
    .B1(_09944_),
    .B2(_09945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_2 _19065_ (.A(_09926_),
    .B(_09955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09956_));
 sky130_fd_sc_hd__a21oi_2 _19066_ (.A1(_09950_),
    .A2(_09952_),
    .B1(_09925_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09957_));
 sky130_fd_sc_hd__nand3_2 _19067_ (.A(_09926_),
    .B(_09954_),
    .C(_09955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09958_));
 sky130_fd_sc_hd__nand3_2 _19068_ (.A(_09925_),
    .B(_09950_),
    .C(_09952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09959_));
 sky130_fd_sc_hd__nand2_2 _19069_ (.A(_09958_),
    .B(_09959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09960_));
 sky130_fd_sc_hd__nand2_2 _19070_ (.A(_09924_),
    .B(_09959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09961_));
 sky130_fd_sc_hd__a21o_2 _19071_ (.A1(_09958_),
    .A2(_09959_),
    .B1(_09924_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09962_));
 sky130_fd_sc_hd__nand2_2 _19072_ (.A(_09837_),
    .B(_09793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09963_));
 sky130_fd_sc_hd__o2bb2ai_2 _19073_ (.A1_N(_09793_),
    .A2_N(_09837_),
    .B1(_09834_),
    .B2(_09828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09964_));
 sky130_fd_sc_hd__o2bb2ai_2 _19074_ (.A1_N(_09794_),
    .A2_N(_09835_),
    .B1(_09836_),
    .B2(_09832_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09965_));
 sky130_fd_sc_hd__o211ai_2 _19075_ (.A1(_09961_),
    .A2(_09957_),
    .B1(_09965_),
    .C1(_09962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09966_));
 sky130_fd_sc_hd__nand4_2 _19076_ (.A(_09922_),
    .B(_09923_),
    .C(_09958_),
    .D(_09959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09967_));
 sky130_fd_sc_hd__a22o_2 _19077_ (.A1(_09922_),
    .A2(_09923_),
    .B1(_09958_),
    .B2(_09959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09968_));
 sky130_fd_sc_hd__a22oi_2 _19078_ (.A1(_09960_),
    .A2(_09924_),
    .B1(_09835_),
    .B2(_09963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09969_));
 sky130_fd_sc_hd__nand3_2 _19079_ (.A(_09968_),
    .B(_09964_),
    .C(_09967_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_2 _19080_ (.A(_09966_),
    .B(_09970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09971_));
 sky130_fd_sc_hd__nand2_2 _19081_ (.A(_09906_),
    .B(_09971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09972_));
 sky130_fd_sc_hd__nand4_2 _19082_ (.A(_09904_),
    .B(_09905_),
    .C(_09966_),
    .D(_09970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09973_));
 sky130_fd_sc_hd__nand3_2 _19083_ (.A(_09906_),
    .B(_09966_),
    .C(_09970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09974_));
 sky130_fd_sc_hd__a21o_2 _19084_ (.A1(_09966_),
    .A2(_09970_),
    .B1(_09906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09975_));
 sky130_fd_sc_hd__nand3_2 _19085_ (.A(_09870_),
    .B(_09974_),
    .C(_09975_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09976_));
 sky130_fd_sc_hd__nand3_2 _19086_ (.A(_09869_),
    .B(_09972_),
    .C(_09973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09977_));
 sky130_fd_sc_hd__a22oi_2 _19087_ (.A1(_09744_),
    .A2(_09745_),
    .B1(_09766_),
    .B2(_09768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09978_));
 sky130_fd_sc_hd__a22o_2 _19088_ (.A1(_09744_),
    .A2(_09745_),
    .B1(_09766_),
    .B2(_09768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09979_));
 sky130_fd_sc_hd__o2111a_2 _19089_ (.A1(_05044_),
    .A2(_06441_),
    .B1(_09745_),
    .C1(_09766_),
    .D1(_09768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09980_));
 sky130_fd_sc_hd__o2111ai_2 _19090_ (.A1(_05044_),
    .A2(_06441_),
    .B1(_09745_),
    .C1(_09766_),
    .D1(_09768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09981_));
 sky130_fd_sc_hd__nor2_2 _19091_ (.A(_09166_),
    .B(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09982_));
 sky130_fd_sc_hd__o22a_2 _19092_ (.A1(_09166_),
    .A2(_09384_),
    .B1(_09978_),
    .B2(_09980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09983_));
 sky130_fd_sc_hd__o22ai_2 _19093_ (.A1(_09166_),
    .A2(_09384_),
    .B1(_09978_),
    .B2(_09980_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09984_));
 sky130_fd_sc_hd__and3_2 _19094_ (.A(_09979_),
    .B(_09981_),
    .C(_09982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09985_));
 sky130_fd_sc_hd__nand4_2 _19095_ (.A(_09979_),
    .B(_09981_),
    .C(\a_l[0] ),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09986_));
 sky130_fd_sc_hd__nand2_2 _19096_ (.A(_09984_),
    .B(_09986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09987_));
 sky130_fd_sc_hd__a21o_2 _19097_ (.A1(_09976_),
    .A2(_09977_),
    .B1(_09987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09988_));
 sky130_fd_sc_hd__o21ai_2 _19098_ (.A1(_09983_),
    .A2(_09985_),
    .B1(_09977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09989_));
 sky130_fd_sc_hd__o211ai_2 _19099_ (.A1(_09983_),
    .A2(_09985_),
    .B1(_09976_),
    .C1(_09977_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09990_));
 sky130_fd_sc_hd__nand3_2 _19100_ (.A(_09868_),
    .B(_09988_),
    .C(_09990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09991_));
 sky130_fd_sc_hd__nand4_2 _19101_ (.A(_09976_),
    .B(_09977_),
    .C(_09984_),
    .D(_09986_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09992_));
 sky130_fd_sc_hd__a21bo_2 _19102_ (.A1(_09976_),
    .A2(_09977_),
    .B1_N(_09987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09993_));
 sky130_fd_sc_hd__a21oi_2 _19103_ (.A1(_09988_),
    .A2(_09990_),
    .B1(_09868_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09994_));
 sky130_fd_sc_hd__nand3_2 _19104_ (.A(_09867_),
    .B(_09992_),
    .C(_09993_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09995_));
 sky130_fd_sc_hd__a21o_2 _19105_ (.A1(_09991_),
    .A2(_09995_),
    .B1(_09736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_09996_));
 sky130_fd_sc_hd__o2111ai_2 _19106_ (.A1(_09625_),
    .A2(_09629_),
    .B1(_09596_),
    .C1(_09991_),
    .D1(_09995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09997_));
 sky130_fd_sc_hd__a21oi_2 _19107_ (.A1(_09996_),
    .A2(_09997_),
    .B1(_09857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09998_));
 sky130_fd_sc_hd__nand3_2 _19108_ (.A(_09996_),
    .B(_09997_),
    .C(_09857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_09999_));
 sky130_fd_sc_hd__nand2b_2 _19109_ (.A_N(_09998_),
    .B(_09999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10000_));
 sky130_fd_sc_hd__a21oi_2 _19110_ (.A1(_09865_),
    .A2(_10000_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10001_));
 sky130_fd_sc_hd__o21a_2 _19111_ (.A1(_09865_),
    .A2(_10000_),
    .B1(_10001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00385_));
 sky130_fd_sc_hd__o21ai_2 _19112_ (.A1(_09860_),
    .A2(_09998_),
    .B1(_09999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10002_));
 sky130_fd_sc_hd__o21a_2 _19113_ (.A1(_09727_),
    .A2(_09859_),
    .B1(_09999_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10003_));
 sky130_fd_sc_hd__nand4_2 _19114_ (.A(_10003_),
    .B(_09734_),
    .C(_09733_),
    .D(_09730_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10004_));
 sky130_fd_sc_hd__nand2_2 _19115_ (.A(_10004_),
    .B(_10002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10005_));
 sky130_fd_sc_hd__a32oi_2 _19116_ (.A1(_09870_),
    .A2(_09974_),
    .A3(_09975_),
    .B1(_09977_),
    .B2(_09987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_2 _19117_ (.A(_09976_),
    .B(_09989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10007_));
 sky130_fd_sc_hd__a22oi_2 _19118_ (.A1(_09969_),
    .A2(_09967_),
    .B1(_09966_),
    .B2(_09906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10008_));
 sky130_fd_sc_hd__o31a_2 _19119_ (.A1(_09253_),
    .A2(_09275_),
    .A3(_04260_),
    .B1(_09915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10009_));
 sky130_fd_sc_hd__a32o_2 _19120_ (.A1(_09910_),
    .A2(\b_l[8] ),
    .A3(\a_l[7] ),
    .B1(_04259_),
    .B2(_06984_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10010_));
 sky130_fd_sc_hd__a21o_2 _19121_ (.A1(_09939_),
    .A2(_09943_),
    .B1(_09940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10011_));
 sky130_fd_sc_hd__a21oi_2 _19122_ (.A1(_09939_),
    .A2(_09943_),
    .B1(_09940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10012_));
 sky130_fd_sc_hd__nand2_2 _19123_ (.A(\a_l[8] ),
    .B(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10013_));
 sky130_fd_sc_hd__nand2_2 _19124_ (.A(\b_l[6] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10014_));
 sky130_fd_sc_hd__nand2_2 _19125_ (.A(\b_l[7] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10015_));
 sky130_fd_sc_hd__a22oi_2 _19126_ (.A1(\b_l[7] ),
    .A2(\a_l[9] ),
    .B1(\a_l[10] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10016_));
 sky130_fd_sc_hd__nand2_2 _19127_ (.A(_10014_),
    .B(_10015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10017_));
 sky130_fd_sc_hd__nand4_2 _19128_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[9] ),
    .D(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10019_));
 sky130_fd_sc_hd__and4_2 _19129_ (.A(_10017_),
    .B(_10019_),
    .C(\a_l[8] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10020_));
 sky130_fd_sc_hd__nand4_2 _19130_ (.A(_10017_),
    .B(_10019_),
    .C(\a_l[8] ),
    .D(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10021_));
 sky130_fd_sc_hd__o2bb2ai_2 _19131_ (.A1_N(_10017_),
    .A2_N(_10019_),
    .B1(_09253_),
    .B2(_09264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10022_));
 sky130_fd_sc_hd__a21o_2 _19132_ (.A1(_10017_),
    .A2(_10019_),
    .B1(_10013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10023_));
 sky130_fd_sc_hd__o211ai_2 _19133_ (.A1(_09253_),
    .A2(_09264_),
    .B1(_10017_),
    .C1(_10019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10024_));
 sky130_fd_sc_hd__nand2_2 _19134_ (.A(_10012_),
    .B(_10022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10025_));
 sky130_fd_sc_hd__nand3_2 _19135_ (.A(_10012_),
    .B(_10021_),
    .C(_10022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10026_));
 sky130_fd_sc_hd__nand3_2 _19136_ (.A(_10023_),
    .B(_10024_),
    .C(_10011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10027_));
 sky130_fd_sc_hd__nand2_2 _19137_ (.A(_10026_),
    .B(_10027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10028_));
 sky130_fd_sc_hd__nand2_2 _19138_ (.A(_10028_),
    .B(_10009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10030_));
 sky130_fd_sc_hd__o211ai_2 _19139_ (.A1(_10020_),
    .A2(_10025_),
    .B1(_10027_),
    .C1(_10010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10031_));
 sky130_fd_sc_hd__nand2_2 _19140_ (.A(_10030_),
    .B(_10031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10032_));
 sky130_fd_sc_hd__o21ai_2 _19141_ (.A1(_09947_),
    .A2(_09948_),
    .B1(_09937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10033_));
 sky130_fd_sc_hd__nand2_2 _19142_ (.A(_09929_),
    .B(_09932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10034_));
 sky130_fd_sc_hd__and4_2 _19143_ (.A(\b_l[1] ),
    .B(\b_l[2] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10035_));
 sky130_fd_sc_hd__nand4_2 _19144_ (.A(\b_l[1] ),
    .B(\b_l[2] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10036_));
 sky130_fd_sc_hd__a22oi_2 _19145_ (.A1(\b_l[2] ),
    .A2(\a_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10037_));
 sky130_fd_sc_hd__a22o_2 _19146_ (.A1(\b_l[2] ),
    .A2(\a_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10038_));
 sky130_fd_sc_hd__nand4_2 _19147_ (.A(_09931_),
    .B(_10034_),
    .C(_10036_),
    .D(_10038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10039_));
 sky130_fd_sc_hd__o2bb2ai_2 _19148_ (.A1_N(_09931_),
    .A2_N(_10034_),
    .B1(_10035_),
    .B2(_10037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10040_));
 sky130_fd_sc_hd__nand2_2 _19149_ (.A(\b_l[5] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10041_));
 sky130_fd_sc_hd__nand2_2 _19150_ (.A(\b_l[3] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10042_));
 sky130_fd_sc_hd__a22oi_2 _19151_ (.A1(\b_l[4] ),
    .A2(\a_l[12] ),
    .B1(\a_l[13] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_2 _19152_ (.A(_09942_),
    .B(_10042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10044_));
 sky130_fd_sc_hd__nand4_2 _19153_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[12] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10045_));
 sky130_fd_sc_hd__a22oi_2 _19154_ (.A1(\b_l[5] ),
    .A2(\a_l[11] ),
    .B1(_10044_),
    .B2(_10045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10046_));
 sky130_fd_sc_hd__and4_2 _19155_ (.A(_10044_),
    .B(_10045_),
    .C(\b_l[5] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10047_));
 sky130_fd_sc_hd__a21oi_2 _19156_ (.A1(_10044_),
    .A2(_10045_),
    .B1(_10041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10048_));
 sky130_fd_sc_hd__a21o_2 _19157_ (.A1(_10044_),
    .A2(_10045_),
    .B1(_10041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10049_));
 sky130_fd_sc_hd__and3_2 _19158_ (.A(_10041_),
    .B(_10044_),
    .C(_10045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10051_));
 sky130_fd_sc_hd__o211ai_2 _19159_ (.A1(_09220_),
    .A2(_09297_),
    .B1(_10044_),
    .C1(_10045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10052_));
 sky130_fd_sc_hd__nand2_2 _19160_ (.A(_10049_),
    .B(_10052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10053_));
 sky130_fd_sc_hd__nand3_2 _19161_ (.A(_10053_),
    .B(_10040_),
    .C(_10039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10054_));
 sky130_fd_sc_hd__o2bb2ai_2 _19162_ (.A1_N(_10039_),
    .A2_N(_10040_),
    .B1(_10046_),
    .B2(_10047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10055_));
 sky130_fd_sc_hd__o211ai_2 _19163_ (.A1(_10046_),
    .A2(_10047_),
    .B1(_10039_),
    .C1(_10040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10056_));
 sky130_fd_sc_hd__o2bb2ai_2 _19164_ (.A1_N(_10039_),
    .A2_N(_10040_),
    .B1(_10048_),
    .B2(_10051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10057_));
 sky130_fd_sc_hd__nand4_2 _19165_ (.A(_09937_),
    .B(_09951_),
    .C(_10054_),
    .D(_10055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10058_));
 sky130_fd_sc_hd__nand4_2 _19166_ (.A(_09938_),
    .B(_10033_),
    .C(_10056_),
    .D(_10057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10059_));
 sky130_fd_sc_hd__nand2_2 _19167_ (.A(_10058_),
    .B(_10059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10060_));
 sky130_fd_sc_hd__nand3_2 _19168_ (.A(_10032_),
    .B(_10058_),
    .C(_10059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10062_));
 sky130_fd_sc_hd__a21o_2 _19169_ (.A1(_10058_),
    .A2(_10059_),
    .B1(_10032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10063_));
 sky130_fd_sc_hd__nand3_2 _19170_ (.A(_10030_),
    .B(_10031_),
    .C(_10059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10064_));
 sky130_fd_sc_hd__nand4_2 _19171_ (.A(_10030_),
    .B(_10031_),
    .C(_10058_),
    .D(_10059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10065_));
 sky130_fd_sc_hd__nand2_2 _19172_ (.A(_10032_),
    .B(_10060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10066_));
 sky130_fd_sc_hd__o2bb2ai_2 _19173_ (.A1_N(_09924_),
    .A2_N(_09959_),
    .B1(_09956_),
    .B2(_09953_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10067_));
 sky130_fd_sc_hd__a21oi_2 _19174_ (.A1(_09924_),
    .A2(_09959_),
    .B1(_09957_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10068_));
 sky130_fd_sc_hd__and3_2 _19175_ (.A(_10067_),
    .B(_10066_),
    .C(_10065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10069_));
 sky130_fd_sc_hd__nand3_2 _19176_ (.A(_10067_),
    .B(_10066_),
    .C(_10065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10070_));
 sky130_fd_sc_hd__nand3_2 _19177_ (.A(_10062_),
    .B(_10063_),
    .C(_10068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10071_));
 sky130_fd_sc_hd__a21oi_2 _19178_ (.A1(_09879_),
    .A2(_09890_),
    .B1(_09893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10073_));
 sky130_fd_sc_hd__a21o_2 _19179_ (.A1(_09879_),
    .A2(_09890_),
    .B1(_09893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10074_));
 sky130_fd_sc_hd__nand2_2 _19180_ (.A(_09918_),
    .B(_09921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10075_));
 sky130_fd_sc_hd__a21boi_2 _19181_ (.A1(_09917_),
    .A2(_09920_),
    .B1_N(_09918_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10076_));
 sky130_fd_sc_hd__nand4_2 _19182_ (.A(\a_l[3] ),
    .B(\a_l[4] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10077_));
 sky130_fd_sc_hd__a22o_2 _19183_ (.A1(\a_l[4] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10078_));
 sky130_fd_sc_hd__and4_2 _19184_ (.A(_10078_),
    .B(\b_l[14] ),
    .C(\a_l[2] ),
    .D(_10077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10079_));
 sky130_fd_sc_hd__o2111ai_2 _19185_ (.A1(_05044_),
    .A2(_06521_),
    .B1(\a_l[2] ),
    .C1(\b_l[14] ),
    .D1(_10078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10080_));
 sky130_fd_sc_hd__o2bb2a_2 _19186_ (.A1_N(_10077_),
    .A2_N(_10078_),
    .B1(_09144_),
    .B2(_09362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10081_));
 sky130_fd_sc_hd__a22o_2 _19187_ (.A1(\a_l[2] ),
    .A2(\b_l[14] ),
    .B1(_10077_),
    .B2(_10078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10082_));
 sky130_fd_sc_hd__nor2_2 _19188_ (.A(_10079_),
    .B(_10081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_2 _19189_ (.A(_10080_),
    .B(_10082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10085_));
 sky130_fd_sc_hd__nand2_2 _19190_ (.A(\a_l[5] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_2 _19191_ (.A(\a_l[6] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_2 _19192_ (.A(\a_l[7] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10088_));
 sky130_fd_sc_hd__nand4_2 _19193_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10089_));
 sky130_fd_sc_hd__a22oi_2 _19194_ (.A1(\a_l[7] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10090_));
 sky130_fd_sc_hd__nand2_2 _19195_ (.A(_10087_),
    .B(_10088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10091_));
 sky130_fd_sc_hd__a21oi_2 _19196_ (.A1(_10089_),
    .A2(_10091_),
    .B1(_10086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10092_));
 sky130_fd_sc_hd__o21ai_2 _19197_ (.A1(_04555_),
    .A2(_06761_),
    .B1(_10086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10093_));
 sky130_fd_sc_hd__o2bb2ai_2 _19198_ (.A1_N(_09885_),
    .A2_N(_09889_),
    .B1(_10090_),
    .B2(_10093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10095_));
 sky130_fd_sc_hd__nand3_2 _19199_ (.A(_10089_),
    .B(\b_l[11] ),
    .C(\a_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10096_));
 sky130_fd_sc_hd__o2bb2ai_2 _19200_ (.A1_N(_10089_),
    .A2_N(_10091_),
    .B1(_09210_),
    .B2(_09308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10097_));
 sky130_fd_sc_hd__o2111ai_2 _19201_ (.A1(_10096_),
    .A2(_10090_),
    .B1(_09889_),
    .C1(_09885_),
    .D1(_10097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10098_));
 sky130_fd_sc_hd__o21ai_2 _19202_ (.A1(_10092_),
    .A2(_10095_),
    .B1(_10098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10099_));
 sky130_fd_sc_hd__o21ai_2 _19203_ (.A1(_10079_),
    .A2(_10081_),
    .B1(_10099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10100_));
 sky130_fd_sc_hd__o2111ai_2 _19204_ (.A1(_10092_),
    .A2(_10095_),
    .B1(_10098_),
    .C1(_10082_),
    .D1(_10080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10101_));
 sky130_fd_sc_hd__o221ai_2 _19205_ (.A1(_10092_),
    .A2(_10095_),
    .B1(_10079_),
    .B2(_10081_),
    .C1(_10098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10102_));
 sky130_fd_sc_hd__nand2_2 _19206_ (.A(_10099_),
    .B(_10084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10103_));
 sky130_fd_sc_hd__nand3_2 _19207_ (.A(_10076_),
    .B(_10102_),
    .C(_10103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10104_));
 sky130_fd_sc_hd__and3_2 _19208_ (.A(_10075_),
    .B(_10100_),
    .C(_10101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10105_));
 sky130_fd_sc_hd__nand3_2 _19209_ (.A(_10075_),
    .B(_10100_),
    .C(_10101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10106_));
 sky130_fd_sc_hd__a31oi_2 _19210_ (.A1(_10076_),
    .A2(_10102_),
    .A3(_10103_),
    .B1(_10073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10107_));
 sky130_fd_sc_hd__a31o_2 _19211_ (.A1(_10076_),
    .A2(_10102_),
    .A3(_10103_),
    .B1(_10073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10108_));
 sky130_fd_sc_hd__a21oi_2 _19212_ (.A1(_10104_),
    .A2(_10106_),
    .B1(_10074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10109_));
 sky130_fd_sc_hd__a21o_2 _19213_ (.A1(_10104_),
    .A2(_10106_),
    .B1(_10074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10110_));
 sky130_fd_sc_hd__and3_2 _19214_ (.A(_10074_),
    .B(_10104_),
    .C(_10106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10111_));
 sky130_fd_sc_hd__nand2_2 _19215_ (.A(_10107_),
    .B(_10106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10112_));
 sky130_fd_sc_hd__o2bb2ai_2 _19216_ (.A1_N(_10070_),
    .A2_N(_10071_),
    .B1(_10109_),
    .B2(_10111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10113_));
 sky130_fd_sc_hd__nand3_2 _19217_ (.A(_10071_),
    .B(_10110_),
    .C(_10112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10114_));
 sky130_fd_sc_hd__nand4_2 _19218_ (.A(_10070_),
    .B(_10071_),
    .C(_10110_),
    .D(_10112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10116_));
 sky130_fd_sc_hd__o211a_2 _19219_ (.A1(_10069_),
    .A2(_10114_),
    .B1(_10113_),
    .C1(_10008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10117_));
 sky130_fd_sc_hd__o211ai_2 _19220_ (.A1(_10069_),
    .A2(_10114_),
    .B1(_10113_),
    .C1(_10008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10118_));
 sky130_fd_sc_hd__a21oi_2 _19221_ (.A1(_10113_),
    .A2(_10116_),
    .B1(_10008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10119_));
 sky130_fd_sc_hd__a21o_2 _19222_ (.A1(_10113_),
    .A2(_10116_),
    .B1(_10008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10120_));
 sky130_fd_sc_hd__nand2_2 _19223_ (.A(\a_l[1] ),
    .B(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10121_));
 sky130_fd_sc_hd__a31o_2 _19224_ (.A1(\a_l[1] ),
    .A2(\b_l[14] ),
    .A3(_09873_),
    .B1(_09874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10122_));
 sky130_fd_sc_hd__o21ai_2 _19225_ (.A1(_09759_),
    .A2(_09902_),
    .B1(_09901_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10123_));
 sky130_fd_sc_hd__o211a_2 _19226_ (.A1(_09874_),
    .A2(_09877_),
    .B1(_09900_),
    .C1(_10123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10124_));
 sky130_fd_sc_hd__o211ai_2 _19227_ (.A1(_09874_),
    .A2(_09877_),
    .B1(_09900_),
    .C1(_10123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10125_));
 sky130_fd_sc_hd__a21oi_2 _19228_ (.A1(_09900_),
    .A2(_10123_),
    .B1(_10122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10127_));
 sky130_fd_sc_hd__o2bb2a_2 _19229_ (.A1_N(\a_l[1] ),
    .A2_N(\b_l[15] ),
    .B1(_10124_),
    .B2(_10127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10128_));
 sky130_fd_sc_hd__o21ai_2 _19230_ (.A1(_10124_),
    .A2(_10127_),
    .B1(_10121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10129_));
 sky130_fd_sc_hd__nor3_2 _19231_ (.A(_10121_),
    .B(_10124_),
    .C(_10127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10130_));
 sky130_fd_sc_hd__nand4b_2 _19232_ (.A_N(_10127_),
    .B(\b_l[15] ),
    .C(\a_l[1] ),
    .D(_10125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10131_));
 sky130_fd_sc_hd__nor2_2 _19233_ (.A(_10128_),
    .B(_10130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10132_));
 sky130_fd_sc_hd__nand2_2 _19234_ (.A(_10129_),
    .B(_10131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10133_));
 sky130_fd_sc_hd__nand2_2 _19235_ (.A(_10132_),
    .B(_10120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10134_));
 sky130_fd_sc_hd__nand4_2 _19236_ (.A(_10118_),
    .B(_10120_),
    .C(_10129_),
    .D(_10131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10135_));
 sky130_fd_sc_hd__o21ai_2 _19237_ (.A1(_10117_),
    .A2(_10119_),
    .B1(_10133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10136_));
 sky130_fd_sc_hd__o21ai_2 _19238_ (.A1(_10117_),
    .A2(_10119_),
    .B1(_10132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10138_));
 sky130_fd_sc_hd__o211ai_2 _19239_ (.A1(_10128_),
    .A2(_10130_),
    .B1(_10118_),
    .C1(_10120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10139_));
 sky130_fd_sc_hd__nand3_2 _19240_ (.A(_10007_),
    .B(_10138_),
    .C(_10139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10140_));
 sky130_fd_sc_hd__nand3_2 _19241_ (.A(_10136_),
    .B(_10006_),
    .C(_10135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10141_));
 sky130_fd_sc_hd__nand2_2 _19242_ (.A(_10140_),
    .B(_10141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10142_));
 sky130_fd_sc_hd__a31o_2 _19243_ (.A1(_09981_),
    .A2(\b_l[15] ),
    .A3(\a_l[0] ),
    .B1(_09978_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10143_));
 sky130_fd_sc_hd__o31a_2 _19244_ (.A1(_09166_),
    .A2(_09384_),
    .A3(_09980_),
    .B1(_09979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10144_));
 sky130_fd_sc_hd__a21o_2 _19245_ (.A1(_10140_),
    .A2(_10141_),
    .B1(_10144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10145_));
 sky130_fd_sc_hd__nand3_2 _19246_ (.A(_10140_),
    .B(_10141_),
    .C(_10144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_2 _19247_ (.A(_10142_),
    .B(_10144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10147_));
 sky130_fd_sc_hd__nand3_2 _19248_ (.A(_10140_),
    .B(_10141_),
    .C(_10143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10149_));
 sky130_fd_sc_hd__a31oi_2 _19249_ (.A1(_09868_),
    .A2(_09988_),
    .A3(_09990_),
    .B1(_09737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10150_));
 sky130_fd_sc_hd__a21oi_2 _19250_ (.A1(_09991_),
    .A2(_09736_),
    .B1(_09994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10151_));
 sky130_fd_sc_hd__nand3_2 _19251_ (.A(_10145_),
    .B(_10146_),
    .C(_10151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10152_));
 sky130_fd_sc_hd__o211ai_2 _19252_ (.A1(_09994_),
    .A2(_10150_),
    .B1(_10149_),
    .C1(_10147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10153_));
 sky130_fd_sc_hd__nand2_2 _19253_ (.A(_10152_),
    .B(_10153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10154_));
 sky130_fd_sc_hd__a21oi_2 _19254_ (.A1(_10005_),
    .A2(_10154_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10155_));
 sky130_fd_sc_hd__o21a_2 _19255_ (.A1(_10005_),
    .A2(_10154_),
    .B1(_10155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00386_));
 sky130_fd_sc_hd__a32oi_2 _19256_ (.A1(_10007_),
    .A2(_10138_),
    .A3(_10139_),
    .B1(_10141_),
    .B2(_10144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10156_));
 sky130_fd_sc_hd__a21boi_2 _19257_ (.A1(_10140_),
    .A2(_10143_),
    .B1_N(_10141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10157_));
 sky130_fd_sc_hd__o21ai_2 _19258_ (.A1(_10133_),
    .A2(_10119_),
    .B1(_10118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10159_));
 sky130_fd_sc_hd__nand2_2 _19259_ (.A(_10058_),
    .B(_10064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10160_));
 sky130_fd_sc_hd__nand3_2 _19260_ (.A(_10039_),
    .B(_10049_),
    .C(_10052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_2 _19261_ (.A(_10040_),
    .B(_10161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10162_));
 sky130_fd_sc_hd__a21o_2 _19262_ (.A1(\b_l[1] ),
    .A2(\a_l[14] ),
    .B1(_09155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10163_));
 sky130_fd_sc_hd__and3_2 _19263_ (.A(_09816_),
    .B(\a_l[15] ),
    .C(\b_l[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10164_));
 sky130_fd_sc_hd__nand2_2 _19264_ (.A(\b_l[5] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10165_));
 sky130_fd_sc_hd__nand2_2 _19265_ (.A(\b_l[4] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10166_));
 sky130_fd_sc_hd__nand2_2 _19266_ (.A(\b_l[3] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10167_));
 sky130_fd_sc_hd__a22o_2 _19267_ (.A1(\b_l[4] ),
    .A2(\a_l[13] ),
    .B1(\a_l[14] ),
    .B2(\b_l[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_10168_));
 sky130_fd_sc_hd__nand2_2 _19268_ (.A(\b_l[4] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10170_));
 sky130_fd_sc_hd__nand4_2 _19269_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[13] ),
    .D(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10171_));
 sky130_fd_sc_hd__o2bb2ai_2 _19270_ (.A1_N(_10166_),
    .A2_N(_10167_),
    .B1(_10170_),
    .B2(_10042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10172_));
 sky130_fd_sc_hd__o221ai_2 _19271_ (.A1(_09220_),
    .A2(_09319_),
    .B1(_10042_),
    .B2(_10170_),
    .C1(_10168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10173_));
 sky130_fd_sc_hd__nand3_2 _19272_ (.A(_10172_),
    .B(\a_l[12] ),
    .C(\b_l[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10174_));
 sky130_fd_sc_hd__nand4_2 _19273_ (.A(_10168_),
    .B(_10171_),
    .C(\b_l[5] ),
    .D(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10175_));
 sky130_fd_sc_hd__o21ai_2 _19274_ (.A1(_09220_),
    .A2(_09319_),
    .B1(_10172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10176_));
 sky130_fd_sc_hd__nand3_2 _19275_ (.A(_10176_),
    .B(_10164_),
    .C(_10175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10177_));
 sky130_fd_sc_hd__o211ai_2 _19276_ (.A1(_09373_),
    .A2(_10163_),
    .B1(_10173_),
    .C1(_10174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_2 _19277_ (.A(_10177_),
    .B(_10178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_10179_));
 sky130_fd_sc_hd__nand4_2 _19278_ (.A(_10040_),
    .B(_10161_),
    .C(_10177_),
    .D(_10178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_2 _19279_ (.A(_10162_),
    .B(_10179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00452_));
 sky130_fd_sc_hd__o21ai_2 _19280_ (.A1(_10041_),
    .A2(_10043_),
    .B1(_10045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00453_));
 sky130_fd_sc_hd__o21a_2 _19281_ (.A1(_10041_),
    .A2(_10043_),
    .B1(_10045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00454_));
 sky130_fd_sc_hd__nand2_2 _19282_ (.A(\b_l[6] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_2 _19283_ (.A(\b_l[7] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00456_));
 sky130_fd_sc_hd__a22oi_2 _19284_ (.A1(\b_l[7] ),
    .A2(\a_l[10] ),
    .B1(\a_l[11] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_2 _19285_ (.A(_00455_),
    .B(_00456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00458_));
 sky130_fd_sc_hd__and3_2 _19286_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(_04259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00459_));
 sky130_fd_sc_hd__nand4_2 _19287_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[10] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_2 _19288_ (.A(\b_l[8] ),
    .B(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00461_));
 sky130_fd_sc_hd__a22o_2 _19289_ (.A1(\b_l[8] ),
    .A2(\a_l[9] ),
    .B1(_00458_),
    .B2(_00460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00462_));
 sky130_fd_sc_hd__and4_2 _19290_ (.A(_00458_),
    .B(_00460_),
    .C(\b_l[8] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00463_));
 sky130_fd_sc_hd__nand4_2 _19291_ (.A(_00458_),
    .B(_00460_),
    .C(\b_l[8] ),
    .D(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00464_));
 sky130_fd_sc_hd__a21o_2 _19292_ (.A1(_00458_),
    .A2(_00460_),
    .B1(_00461_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00465_));
 sky130_fd_sc_hd__o211ai_2 _19293_ (.A1(_09264_),
    .A2(_09275_),
    .B1(_00458_),
    .C1(_00460_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00466_));
 sky130_fd_sc_hd__nand3_2 _19294_ (.A(_00454_),
    .B(_00465_),
    .C(_00466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_2 _19295_ (.A(_00462_),
    .B(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00468_));
 sky130_fd_sc_hd__nand3_2 _19296_ (.A(_00462_),
    .B(_00464_),
    .C(_00453_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00469_));
 sky130_fd_sc_hd__o21ai_2 _19297_ (.A1(_10013_),
    .A2(_10016_),
    .B1(_10019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00470_));
 sky130_fd_sc_hd__a21boi_2 _19298_ (.A1(_00467_),
    .A2(_00469_),
    .B1_N(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00472_));
 sky130_fd_sc_hd__a21bo_2 _19299_ (.A1(_00467_),
    .A2(_00469_),
    .B1_N(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00473_));
 sky130_fd_sc_hd__o2111a_2 _19300_ (.A1(_10013_),
    .A2(_10016_),
    .B1(_10019_),
    .C1(_00467_),
    .D1(_00469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00474_));
 sky130_fd_sc_hd__o2111ai_2 _19301_ (.A1(_10013_),
    .A2(_10016_),
    .B1(_10019_),
    .C1(_00467_),
    .D1(_00469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00475_));
 sky130_fd_sc_hd__a21oi_2 _19302_ (.A1(_00467_),
    .A2(_00469_),
    .B1(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00476_));
 sky130_fd_sc_hd__a21o_2 _19303_ (.A1(_00467_),
    .A2(_00469_),
    .B1(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00477_));
 sky130_fd_sc_hd__and3_2 _19304_ (.A(_00467_),
    .B(_00469_),
    .C(_00470_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00478_));
 sky130_fd_sc_hd__o211ai_2 _19305_ (.A1(_00463_),
    .A2(_00468_),
    .B1(_00470_),
    .C1(_00467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00479_));
 sky130_fd_sc_hd__nand4_2 _19306_ (.A(_00451_),
    .B(_00452_),
    .C(_00477_),
    .D(_00479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00480_));
 sky130_fd_sc_hd__o2bb2ai_2 _19307_ (.A1_N(_00451_),
    .A2_N(_00452_),
    .B1(_00476_),
    .B2(_00478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00481_));
 sky130_fd_sc_hd__o2bb2ai_2 _19308_ (.A1_N(_00451_),
    .A2_N(_00452_),
    .B1(_00472_),
    .B2(_00474_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00483_));
 sky130_fd_sc_hd__o211ai_2 _19309_ (.A1(_10179_),
    .A2(_10162_),
    .B1(_00475_),
    .C1(_00473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00484_));
 sky130_fd_sc_hd__nand4_2 _19310_ (.A(_00451_),
    .B(_00452_),
    .C(_00473_),
    .D(_00475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_2 _19311_ (.A(_00483_),
    .B(_00485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_2 _19312_ (.A(_10032_),
    .B(_10058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00487_));
 sky130_fd_sc_hd__nand4_2 _19313_ (.A(_10059_),
    .B(_00480_),
    .C(_00481_),
    .D(_00487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00488_));
 sky130_fd_sc_hd__and4_2 _19314_ (.A(_10058_),
    .B(_10064_),
    .C(_00483_),
    .D(_00485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00489_));
 sky130_fd_sc_hd__nand4_2 _19315_ (.A(_10058_),
    .B(_10064_),
    .C(_00483_),
    .D(_00485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00490_));
 sky130_fd_sc_hd__nand2_2 _19316_ (.A(_00488_),
    .B(_00490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00491_));
 sky130_fd_sc_hd__o2bb2ai_2 _19317_ (.A1_N(_10010_),
    .A2_N(_10027_),
    .B1(_10025_),
    .B2(_10020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00492_));
 sky130_fd_sc_hd__a21boi_2 _19318_ (.A1(_10010_),
    .A2(_10027_),
    .B1_N(_10026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00494_));
 sky130_fd_sc_hd__a21o_2 _19319_ (.A1(_10086_),
    .A2(_10089_),
    .B1(_10090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00495_));
 sky130_fd_sc_hd__nand2_2 _19320_ (.A(\a_l[6] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_2 _19321_ (.A(\a_l[7] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_2 _19322_ (.A(\a_l[8] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00498_));
 sky130_fd_sc_hd__a22oi_2 _19323_ (.A1(\a_l[8] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_2 _19324_ (.A(_00497_),
    .B(_00498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00500_));
 sky130_fd_sc_hd__nand4_2 _19325_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00501_));
 sky130_fd_sc_hd__a21o_2 _19326_ (.A1(_00500_),
    .A2(_00501_),
    .B1(_00496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00502_));
 sky130_fd_sc_hd__o211ai_2 _19327_ (.A1(_09231_),
    .A2(_09308_),
    .B1(_00500_),
    .C1(_00501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00503_));
 sky130_fd_sc_hd__a22oi_2 _19328_ (.A1(\a_l[6] ),
    .A2(\b_l[11] ),
    .B1(_00500_),
    .B2(_00501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00505_));
 sky130_fd_sc_hd__nand3_2 _19329_ (.A(_00501_),
    .B(\b_l[11] ),
    .C(\a_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00506_));
 sky130_fd_sc_hd__nand3_2 _19330_ (.A(_00502_),
    .B(_00503_),
    .C(_00495_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00507_));
 sky130_fd_sc_hd__and3_2 _19331_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00508_));
 sky130_fd_sc_hd__nand4_2 _19332_ (.A(\a_l[4] ),
    .B(\a_l[5] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00509_));
 sky130_fd_sc_hd__a22o_2 _19333_ (.A1(\a_l[5] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00510_));
 sky130_fd_sc_hd__o2111a_2 _19334_ (.A1(_05044_),
    .A2(_06605_),
    .B1(\a_l[3] ),
    .C1(\b_l[14] ),
    .D1(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00511_));
 sky130_fd_sc_hd__o2111ai_2 _19335_ (.A1(_05044_),
    .A2(_06605_),
    .B1(\a_l[3] ),
    .C1(\b_l[14] ),
    .D1(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00512_));
 sky130_fd_sc_hd__a22oi_2 _19336_ (.A1(\a_l[3] ),
    .A2(\b_l[14] ),
    .B1(_00509_),
    .B2(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00513_));
 sky130_fd_sc_hd__a22o_2 _19337_ (.A1(\a_l[3] ),
    .A2(\b_l[14] ),
    .B1(_00509_),
    .B2(_00510_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00514_));
 sky130_fd_sc_hd__nor2_2 _19338_ (.A(_00511_),
    .B(_00513_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_2 _19339_ (.A(_00512_),
    .B(_00514_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00517_));
 sky130_fd_sc_hd__o211ai_2 _19340_ (.A1(_00499_),
    .A2(_00506_),
    .B1(_10091_),
    .C1(_10093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00518_));
 sky130_fd_sc_hd__o21ai_2 _19341_ (.A1(_00505_),
    .A2(_00518_),
    .B1(_00507_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00519_));
 sky130_fd_sc_hd__o211ai_2 _19342_ (.A1(_00518_),
    .A2(_00505_),
    .B1(_00507_),
    .C1(_00517_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_2 _19343_ (.A(_00519_),
    .B(_00516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00521_));
 sky130_fd_sc_hd__o21ai_2 _19344_ (.A1(_00511_),
    .A2(_00513_),
    .B1(_00519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00522_));
 sky130_fd_sc_hd__o211ai_2 _19345_ (.A1(_00505_),
    .A2(_00518_),
    .B1(_00507_),
    .C1(_00516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00523_));
 sky130_fd_sc_hd__nand3_2 _19346_ (.A(_00494_),
    .B(_00520_),
    .C(_00521_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00524_));
 sky130_fd_sc_hd__nand3_2 _19347_ (.A(_00522_),
    .B(_00523_),
    .C(_00492_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00525_));
 sky130_fd_sc_hd__o2bb2a_2 _19348_ (.A1_N(_10085_),
    .A2_N(_10098_),
    .B1(_10095_),
    .B2(_10092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00526_));
 sky130_fd_sc_hd__a2bb2o_2 _19349_ (.A1_N(_10092_),
    .A2_N(_10095_),
    .B1(_10098_),
    .B2(_10085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00527_));
 sky130_fd_sc_hd__a21o_2 _19350_ (.A1(_00524_),
    .A2(_00525_),
    .B1(_00526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00528_));
 sky130_fd_sc_hd__nand3_2 _19351_ (.A(_00524_),
    .B(_00525_),
    .C(_00526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00529_));
 sky130_fd_sc_hd__a21o_2 _19352_ (.A1(_00524_),
    .A2(_00525_),
    .B1(_00527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00530_));
 sky130_fd_sc_hd__nand3_2 _19353_ (.A(_00524_),
    .B(_00525_),
    .C(_00527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_2 _19354_ (.A(_00530_),
    .B(_00531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_2 _19355_ (.A(_00528_),
    .B(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_2 _19356_ (.A(_00491_),
    .B(_00532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00534_));
 sky130_fd_sc_hd__nand4_2 _19357_ (.A(_00488_),
    .B(_00490_),
    .C(_00530_),
    .D(_00531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00535_));
 sky130_fd_sc_hd__a21oi_2 _19358_ (.A1(_00488_),
    .A2(_00490_),
    .B1(_00532_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00537_));
 sky130_fd_sc_hd__nand2_2 _19359_ (.A(_00491_),
    .B(_00533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00538_));
 sky130_fd_sc_hd__nand4_2 _19360_ (.A(_00488_),
    .B(_00490_),
    .C(_00528_),
    .D(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00539_));
 sky130_fd_sc_hd__o21ai_2 _19361_ (.A1(_10109_),
    .A2(_10111_),
    .B1(_10070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00540_));
 sky130_fd_sc_hd__a22oi_2 _19362_ (.A1(_00538_),
    .A2(_00539_),
    .B1(_00540_),
    .B2(_10071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00541_));
 sky130_fd_sc_hd__nand4_2 _19363_ (.A(_10070_),
    .B(_10114_),
    .C(_00534_),
    .D(_00535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00542_));
 sky130_fd_sc_hd__nand3_2 _19364_ (.A(_10071_),
    .B(_00539_),
    .C(_00540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00543_));
 sky130_fd_sc_hd__nand4_2 _19365_ (.A(_10071_),
    .B(_00538_),
    .C(_00539_),
    .D(_00540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_2 _19366_ (.A(_09144_),
    .B(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00545_));
 sky130_fd_sc_hd__o2bb2ai_2 _19367_ (.A1_N(_10077_),
    .A2_N(_10080_),
    .B1(_10105_),
    .B2(_10107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00546_));
 sky130_fd_sc_hd__o2111ai_2 _19368_ (.A1(_05044_),
    .A2(_06521_),
    .B1(_10080_),
    .C1(_10106_),
    .D1(_10108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _19369_ (.A(_00548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00549_));
 sky130_fd_sc_hd__a21oi_2 _19370_ (.A1(_00546_),
    .A2(_00548_),
    .B1(_00545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00550_));
 sky130_fd_sc_hd__a22o_2 _19371_ (.A1(\a_l[2] ),
    .A2(\b_l[15] ),
    .B1(_00546_),
    .B2(_00548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00551_));
 sky130_fd_sc_hd__and3_2 _19372_ (.A(_00546_),
    .B(_00548_),
    .C(_00545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00552_));
 sky130_fd_sc_hd__nand4_2 _19373_ (.A(_00546_),
    .B(_00548_),
    .C(\a_l[2] ),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00553_));
 sky130_fd_sc_hd__nor2_2 _19374_ (.A(_00550_),
    .B(_00552_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_2 _19375_ (.A(_00551_),
    .B(_00553_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00555_));
 sky130_fd_sc_hd__a21o_2 _19376_ (.A1(_00542_),
    .A2(_00544_),
    .B1(_00555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00556_));
 sky130_fd_sc_hd__o211ai_2 _19377_ (.A1(_00537_),
    .A2(_00543_),
    .B1(_00555_),
    .C1(_00542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00557_));
 sky130_fd_sc_hd__o2111ai_2 _19378_ (.A1(_00537_),
    .A2(_00543_),
    .B1(_00551_),
    .C1(_00553_),
    .D1(_00542_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00559_));
 sky130_fd_sc_hd__a21o_2 _19379_ (.A1(_00542_),
    .A2(_00544_),
    .B1(_00554_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00560_));
 sky130_fd_sc_hd__nand4_2 _19380_ (.A(_10118_),
    .B(_10134_),
    .C(_00556_),
    .D(_00557_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00561_));
 sky130_fd_sc_hd__nand3_2 _19381_ (.A(_00560_),
    .B(_10159_),
    .C(_00559_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00562_));
 sky130_fd_sc_hd__o21ai_2 _19382_ (.A1(_10121_),
    .A2(_10127_),
    .B1(_10125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00563_));
 sky130_fd_sc_hd__o21a_2 _19383_ (.A1(_10121_),
    .A2(_10127_),
    .B1(_10125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00564_));
 sky130_fd_sc_hd__a21o_2 _19384_ (.A1(_00561_),
    .A2(_00562_),
    .B1(_00563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00565_));
 sky130_fd_sc_hd__nand3_2 _19385_ (.A(_00561_),
    .B(_00562_),
    .C(_00563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00566_));
 sky130_fd_sc_hd__o2111ai_2 _19386_ (.A1(_10127_),
    .A2(_10121_),
    .B1(_10125_),
    .C1(_00561_),
    .D1(_00562_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00567_));
 sky130_fd_sc_hd__a21o_2 _19387_ (.A1(_00561_),
    .A2(_00562_),
    .B1(_00564_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00568_));
 sky130_fd_sc_hd__nand3_2 _19388_ (.A(_10157_),
    .B(_00567_),
    .C(_00568_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00570_));
 sky130_fd_sc_hd__nand3_2 _19389_ (.A(_10156_),
    .B(_00565_),
    .C(_00566_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_2 _19390_ (.A(_00570_),
    .B(_00571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_2 _19391_ (.A(_10005_),
    .B(_10153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_2 _19392_ (.A(_10152_),
    .B(_00573_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00574_));
 sky130_fd_sc_hd__a21oi_2 _19393_ (.A1(_00572_),
    .A2(_00574_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00575_));
 sky130_fd_sc_hd__o21a_2 _19394_ (.A1(_00572_),
    .A2(_00574_),
    .B1(_00575_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00387_));
 sky130_fd_sc_hd__a31o_2 _19395_ (.A1(_00560_),
    .A2(_10159_),
    .A3(_00559_),
    .B1(_00563_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00576_));
 sky130_fd_sc_hd__o22ai_2 _19396_ (.A1(_00537_),
    .A2(_00543_),
    .B1(_00555_),
    .B2(_00541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00577_));
 sky130_fd_sc_hd__a21boi_2 _19397_ (.A1(_00554_),
    .A2(_00542_),
    .B1_N(_00544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00578_));
 sky130_fd_sc_hd__nor2_2 _19398_ (.A(_09188_),
    .B(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_2 _19399_ (.A(_00525_),
    .B(_00527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_2 _19400_ (.A(_00524_),
    .B(_00526_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00582_));
 sky130_fd_sc_hd__o211ai_2 _19401_ (.A1(_00508_),
    .A2(_00511_),
    .B1(_00524_),
    .C1(_00581_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00583_));
 sky130_fd_sc_hd__inv_2 _19402_ (.A(_00583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00584_));
 sky130_fd_sc_hd__o2111ai_2 _19403_ (.A1(_05044_),
    .A2(_06605_),
    .B1(_00512_),
    .C1(_00525_),
    .D1(_00582_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00585_));
 sky130_fd_sc_hd__a21oi_2 _19404_ (.A1(_00583_),
    .A2(_00585_),
    .B1(_00580_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00586_));
 sky130_fd_sc_hd__and3_2 _19405_ (.A(_00585_),
    .B(_00580_),
    .C(_00583_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00587_));
 sky130_fd_sc_hd__nor2_2 _19406_ (.A(_00586_),
    .B(_00587_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00588_));
 sky130_fd_sc_hd__a2bb2o_2 _19407_ (.A1_N(_00505_),
    .A2_N(_00518_),
    .B1(_00507_),
    .B2(_00516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00589_));
 sky130_fd_sc_hd__o2bb2ai_2 _19408_ (.A1_N(_00470_),
    .A2_N(_00467_),
    .B1(_00463_),
    .B2(_00468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00591_));
 sky130_fd_sc_hd__a21boi_2 _19409_ (.A1(_00467_),
    .A2(_00470_),
    .B1_N(_00469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00592_));
 sky130_fd_sc_hd__a21o_2 _19410_ (.A1(_00496_),
    .A2(_00501_),
    .B1(_00499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00593_));
 sky130_fd_sc_hd__a21oi_2 _19411_ (.A1(_00496_),
    .A2(_00501_),
    .B1(_00499_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_2 _19412_ (.A(\a_l[7] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_2 _19413_ (.A(\a_l[8] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_2 _19414_ (.A(\a_l[9] ),
    .B(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00597_));
 sky130_fd_sc_hd__a22oi_2 _19415_ (.A1(\a_l[9] ),
    .A2(\b_l[9] ),
    .B1(\b_l[10] ),
    .B2(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_2 _19416_ (.A(_00596_),
    .B(_00597_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00599_));
 sky130_fd_sc_hd__nor2_2 _19417_ (.A(_04555_),
    .B(_06985_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00600_));
 sky130_fd_sc_hd__nand4_2 _19418_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .C(\b_l[9] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00601_));
 sky130_fd_sc_hd__a41o_2 _19419_ (.A1(\a_l[8] ),
    .A2(\a_l[9] ),
    .A3(\b_l[9] ),
    .A4(\b_l[10] ),
    .B1(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00602_));
 sky130_fd_sc_hd__o21ai_2 _19420_ (.A1(_00598_),
    .A2(_00600_),
    .B1(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00603_));
 sky130_fd_sc_hd__o221ai_2 _19421_ (.A1(_09242_),
    .A2(_09308_),
    .B1(_04555_),
    .B2(_06985_),
    .C1(_00599_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00604_));
 sky130_fd_sc_hd__a21o_2 _19422_ (.A1(_00599_),
    .A2(_00601_),
    .B1(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00605_));
 sky130_fd_sc_hd__o211a_2 _19423_ (.A1(_00602_),
    .A2(_00598_),
    .B1(_00594_),
    .C1(_00603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00606_));
 sky130_fd_sc_hd__o211ai_2 _19424_ (.A1(_00602_),
    .A2(_00598_),
    .B1(_00594_),
    .C1(_00603_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00607_));
 sky130_fd_sc_hd__nand3_2 _19425_ (.A(_00605_),
    .B(_00593_),
    .C(_00604_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00608_));
 sky130_fd_sc_hd__inv_2 _19426_ (.A(_00608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_2 _19427_ (.A(\a_l[4] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_2 _19428_ (.A(\a_l[5] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_2 _19429_ (.A(\a_l[6] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00613_));
 sky130_fd_sc_hd__nand4_2 _19430_ (.A(\a_l[5] ),
    .B(\a_l[6] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00614_));
 sky130_fd_sc_hd__o22a_2 _19431_ (.A1(_09231_),
    .A2(_09329_),
    .B1(_09351_),
    .B2(_09210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00615_));
 sky130_fd_sc_hd__nand2_2 _19432_ (.A(_00612_),
    .B(_00613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00616_));
 sky130_fd_sc_hd__o2bb2a_2 _19433_ (.A1_N(_00614_),
    .A2_N(_00616_),
    .B1(_09199_),
    .B2(_09362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00617_));
 sky130_fd_sc_hd__and4_2 _19434_ (.A(_00616_),
    .B(\b_l[14] ),
    .C(\a_l[4] ),
    .D(_00614_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00618_));
 sky130_fd_sc_hd__a21oi_2 _19435_ (.A1(_00614_),
    .A2(_00616_),
    .B1(_00610_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00619_));
 sky130_fd_sc_hd__o22a_2 _19436_ (.A1(_09199_),
    .A2(_09362_),
    .B1(_00612_),
    .B2(_00613_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00620_));
 sky130_fd_sc_hd__a21o_2 _19437_ (.A1(_00616_),
    .A2(_00620_),
    .B1(_00619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00621_));
 sky130_fd_sc_hd__a21oi_2 _19438_ (.A1(_00620_),
    .A2(_00616_),
    .B1(_00619_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00623_));
 sky130_fd_sc_hd__a21o_2 _19439_ (.A1(_00607_),
    .A2(_00608_),
    .B1(_00623_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00624_));
 sky130_fd_sc_hd__o211ai_2 _19440_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_00607_),
    .C1(_00608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00625_));
 sky130_fd_sc_hd__o2bb2ai_2 _19441_ (.A1_N(_00607_),
    .A2_N(_00608_),
    .B1(_00617_),
    .B2(_00618_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00626_));
 sky130_fd_sc_hd__nand3_2 _19442_ (.A(_00621_),
    .B(_00608_),
    .C(_00607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00627_));
 sky130_fd_sc_hd__nand3_2 _19443_ (.A(_00592_),
    .B(_00624_),
    .C(_00625_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00628_));
 sky130_fd_sc_hd__a21oi_2 _19444_ (.A1(_00624_),
    .A2(_00625_),
    .B1(_00592_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00629_));
 sky130_fd_sc_hd__nand3_2 _19445_ (.A(_00626_),
    .B(_00627_),
    .C(_00591_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00630_));
 sky130_fd_sc_hd__a21o_2 _19446_ (.A1(_00628_),
    .A2(_00630_),
    .B1(_00589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00631_));
 sky130_fd_sc_hd__nand2_2 _19447_ (.A(_00628_),
    .B(_00589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00632_));
 sky130_fd_sc_hd__nand3_2 _19448_ (.A(_00628_),
    .B(_00630_),
    .C(_00589_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00634_));
 sky130_fd_sc_hd__o21ai_2 _19449_ (.A1(_00629_),
    .A2(_00632_),
    .B1(_00631_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_2 _19450_ (.A(\b_l[5] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_2 _19451_ (.A(\b_l[3] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_2 _19452_ (.A(_10170_),
    .B(_00637_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00638_));
 sky130_fd_sc_hd__nand4_2 _19453_ (.A(\b_l[3] ),
    .B(\b_l[4] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00639_));
 sky130_fd_sc_hd__and3_2 _19454_ (.A(_00636_),
    .B(_00638_),
    .C(_00639_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00640_));
 sky130_fd_sc_hd__a21oi_2 _19455_ (.A1(_00638_),
    .A2(_00639_),
    .B1(_00636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00641_));
 sky130_fd_sc_hd__nor2_2 _19456_ (.A(_00640_),
    .B(_00641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00642_));
 sky130_fd_sc_hd__o2bb2ai_2 _19457_ (.A1_N(_10036_),
    .A2_N(_10177_),
    .B1(_00640_),
    .B2(_00641_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00643_));
 sky130_fd_sc_hd__nand3_2 _19458_ (.A(_00642_),
    .B(_10177_),
    .C(_10036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00645_));
 sky130_fd_sc_hd__inv_2 _19459_ (.A(_00645_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00646_));
 sky130_fd_sc_hd__a22oi_2 _19460_ (.A1(_10166_),
    .A2(_10167_),
    .B1(_10171_),
    .B2(_10165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00647_));
 sky130_fd_sc_hd__a22o_2 _19461_ (.A1(_10166_),
    .A2(_10167_),
    .B1(_10171_),
    .B2(_10165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00648_));
 sky130_fd_sc_hd__nand2_2 _19462_ (.A(\b_l[6] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_2 _19463_ (.A(\b_l[7] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00650_));
 sky130_fd_sc_hd__a22oi_2 _19464_ (.A1(\b_l[7] ),
    .A2(\a_l[11] ),
    .B1(\a_l[12] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00651_));
 sky130_fd_sc_hd__a22o_2 _19465_ (.A1(\b_l[7] ),
    .A2(\a_l[11] ),
    .B1(\a_l[12] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00652_));
 sky130_fd_sc_hd__nand2_2 _19466_ (.A(\b_l[7] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00653_));
 sky130_fd_sc_hd__o2bb2ai_2 _19467_ (.A1_N(_00649_),
    .A2_N(_00650_),
    .B1(_00653_),
    .B2(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00654_));
 sky130_fd_sc_hd__and2_2 _19468_ (.A(\b_l[8] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00656_));
 sky130_fd_sc_hd__o21ai_2 _19469_ (.A1(_09264_),
    .A2(_09286_),
    .B1(_00654_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00657_));
 sky130_fd_sc_hd__o211ai_2 _19470_ (.A1(_00455_),
    .A2(_00653_),
    .B1(_00656_),
    .C1(_00652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00658_));
 sky130_fd_sc_hd__o221ai_2 _19471_ (.A1(_09264_),
    .A2(_09286_),
    .B1(_00455_),
    .B2(_00653_),
    .C1(_00652_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_2 _19472_ (.A(_00654_),
    .B(_00656_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00660_));
 sky130_fd_sc_hd__nand3_2 _19473_ (.A(_00648_),
    .B(_00659_),
    .C(_00660_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00661_));
 sky130_fd_sc_hd__nand3_2 _19474_ (.A(_00657_),
    .B(_00658_),
    .C(_00647_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00662_));
 sky130_fd_sc_hd__and3_2 _19475_ (.A(_00458_),
    .B(\a_l[9] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00663_));
 sky130_fd_sc_hd__a21o_2 _19476_ (.A1(_00460_),
    .A2(_00461_),
    .B1(_00457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00664_));
 sky130_fd_sc_hd__a21oi_2 _19477_ (.A1(_00460_),
    .A2(_00461_),
    .B1(_00457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00665_));
 sky130_fd_sc_hd__a21oi_2 _19478_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00666_));
 sky130_fd_sc_hd__a21o_2 _19479_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00667_));
 sky130_fd_sc_hd__and3_2 _19480_ (.A(_00661_),
    .B(_00662_),
    .C(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00668_));
 sky130_fd_sc_hd__nand3_2 _19481_ (.A(_00661_),
    .B(_00662_),
    .C(_00664_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00669_));
 sky130_fd_sc_hd__a21oi_2 _19482_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00670_));
 sky130_fd_sc_hd__a21o_2 _19483_ (.A1(_00661_),
    .A2(_00662_),
    .B1(_00665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00671_));
 sky130_fd_sc_hd__and3_2 _19484_ (.A(_00661_),
    .B(_00662_),
    .C(_00665_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00672_));
 sky130_fd_sc_hd__o211ai_2 _19485_ (.A1(_00459_),
    .A2(_00663_),
    .B1(_00662_),
    .C1(_00661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00673_));
 sky130_fd_sc_hd__o2bb2ai_2 _19486_ (.A1_N(_00643_),
    .A2_N(_00645_),
    .B1(_00670_),
    .B2(_00672_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00674_));
 sky130_fd_sc_hd__nand4_2 _19487_ (.A(_00643_),
    .B(_00645_),
    .C(_00671_),
    .D(_00673_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00675_));
 sky130_fd_sc_hd__o2bb2ai_2 _19488_ (.A1_N(_00643_),
    .A2_N(_00645_),
    .B1(_00666_),
    .B2(_00668_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00677_));
 sky130_fd_sc_hd__nand4_2 _19489_ (.A(_00643_),
    .B(_00645_),
    .C(_00667_),
    .D(_00669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00678_));
 sky130_fd_sc_hd__nand3_2 _19490_ (.A(_00452_),
    .B(_00477_),
    .C(_00479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00679_));
 sky130_fd_sc_hd__a22oi_2 _19491_ (.A1(_00677_),
    .A2(_00678_),
    .B1(_00679_),
    .B2(_00451_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00680_));
 sky130_fd_sc_hd__nand4_2 _19492_ (.A(_00452_),
    .B(_00484_),
    .C(_00674_),
    .D(_00675_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00681_));
 sky130_fd_sc_hd__nand4_2 _19493_ (.A(_00451_),
    .B(_00677_),
    .C(_00678_),
    .D(_00679_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_2 _19494_ (.A(_00681_),
    .B(_00682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00683_));
 sky130_fd_sc_hd__nand4_2 _19495_ (.A(_00631_),
    .B(_00634_),
    .C(_00681_),
    .D(_00682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00684_));
 sky130_fd_sc_hd__a22oi_2 _19496_ (.A1(_00631_),
    .A2(_00634_),
    .B1(_00681_),
    .B2(_00682_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_2 _19497_ (.A(_00635_),
    .B(_00683_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3_2 _19498_ (.A(_00490_),
    .B(_00528_),
    .C(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00688_));
 sky130_fd_sc_hd__a22oi_2 _19499_ (.A1(_10160_),
    .A2(_00486_),
    .B1(_00528_),
    .B2(_00529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00689_));
 sky130_fd_sc_hd__nand3_2 _19500_ (.A(_00488_),
    .B(_00530_),
    .C(_00531_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00690_));
 sky130_fd_sc_hd__nand2_2 _19501_ (.A(_00488_),
    .B(_00688_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00691_));
 sky130_fd_sc_hd__a21oi_2 _19502_ (.A1(_00684_),
    .A2(_00686_),
    .B1(_00691_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00692_));
 sky130_fd_sc_hd__o2bb2ai_2 _19503_ (.A1_N(_00684_),
    .A2_N(_00686_),
    .B1(_00689_),
    .B2(_00489_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00693_));
 sky130_fd_sc_hd__o211ai_2 _19504_ (.A1(_00486_),
    .A2(_10160_),
    .B1(_00690_),
    .C1(_00684_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00694_));
 sky130_fd_sc_hd__nor2_2 _19505_ (.A(_00685_),
    .B(_00694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00695_));
 sky130_fd_sc_hd__o22ai_2 _19506_ (.A1(_00586_),
    .A2(_00587_),
    .B1(_00692_),
    .B2(_00695_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_2 _19507_ (.A(_00693_),
    .B(_00588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00697_));
 sky130_fd_sc_hd__o221ai_2 _19508_ (.A1(_00586_),
    .A2(_00587_),
    .B1(_00685_),
    .B2(_00694_),
    .C1(_00693_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00699_));
 sky130_fd_sc_hd__o21ai_2 _19509_ (.A1(_00692_),
    .A2(_00695_),
    .B1(_00588_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00700_));
 sky130_fd_sc_hd__o211ai_2 _19510_ (.A1(_00695_),
    .A2(_00697_),
    .B1(_00696_),
    .C1(_00577_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00701_));
 sky130_fd_sc_hd__nand3_2 _19511_ (.A(_00578_),
    .B(_00699_),
    .C(_00700_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00702_));
 sky130_fd_sc_hd__o21a_2 _19512_ (.A1(_09144_),
    .A2(_09384_),
    .B1(_00546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00703_));
 sky130_fd_sc_hd__o21ai_2 _19513_ (.A1(_09144_),
    .A2(_09384_),
    .B1(_00546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00704_));
 sky130_fd_sc_hd__o2bb2ai_2 _19514_ (.A1_N(_00701_),
    .A2_N(_00702_),
    .B1(_00703_),
    .B2(_00549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00705_));
 sky130_fd_sc_hd__nand4_2 _19515_ (.A(_00548_),
    .B(_00701_),
    .C(_00702_),
    .D(_00704_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00706_));
 sky130_fd_sc_hd__a22o_2 _19516_ (.A1(_00561_),
    .A2(_00576_),
    .B1(_00705_),
    .B2(_00706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00707_));
 sky130_fd_sc_hd__nand4_2 _19517_ (.A(_00561_),
    .B(_00576_),
    .C(_00705_),
    .D(_00706_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_2 _19518_ (.A(_00707_),
    .B(_00708_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00710_));
 sky130_fd_sc_hd__and4_2 _19519_ (.A(_10152_),
    .B(_10153_),
    .C(_00570_),
    .D(_00571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00711_));
 sky130_fd_sc_hd__nand4_2 _19520_ (.A(_10152_),
    .B(_10153_),
    .C(_00570_),
    .D(_00571_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00712_));
 sky130_fd_sc_hd__a21boi_2 _19521_ (.A1(_10153_),
    .A2(_00571_),
    .B1_N(_00570_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00713_));
 sky130_fd_sc_hd__a31o_2 _19522_ (.A1(_10004_),
    .A2(_00711_),
    .A3(_10002_),
    .B1(_00713_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00714_));
 sky130_fd_sc_hd__a21oi_2 _19523_ (.A1(_00707_),
    .A2(_00708_),
    .B1(_00714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00715_));
 sky130_fd_sc_hd__nand3_2 _19524_ (.A(_00707_),
    .B(_00708_),
    .C(_00714_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00716_));
 sky130_fd_sc_hd__nor3b_2 _19525_ (.A(rst),
    .B(_00715_),
    .C_N(_00716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00388_));
 sky130_fd_sc_hd__a21oi_2 _19526_ (.A1(_00580_),
    .A2(_00585_),
    .B1(_00584_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00717_));
 sky130_fd_sc_hd__o22ai_2 _19527_ (.A1(_00586_),
    .A2(_00587_),
    .B1(_00685_),
    .B2(_00694_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_2 _19528_ (.A(_00693_),
    .B(_00718_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00720_));
 sky130_fd_sc_hd__o21ai_2 _19529_ (.A1(_00685_),
    .A2(_00694_),
    .B1(_00697_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00721_));
 sky130_fd_sc_hd__nand2_2 _19530_ (.A(\a_l[4] ),
    .B(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00722_));
 sky130_fd_sc_hd__a21oi_2 _19531_ (.A1(_00610_),
    .A2(_00614_),
    .B1(_00615_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00723_));
 sky130_fd_sc_hd__o211ai_2 _19532_ (.A1(_00589_),
    .A2(_00629_),
    .B1(_00723_),
    .C1(_00628_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00724_));
 sky130_fd_sc_hd__o211ai_2 _19533_ (.A1(_00615_),
    .A2(_00620_),
    .B1(_00630_),
    .C1(_00632_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00725_));
 sky130_fd_sc_hd__a21o_2 _19534_ (.A1(_00724_),
    .A2(_00725_),
    .B1(_00722_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00726_));
 sky130_fd_sc_hd__o21ai_2 _19535_ (.A1(_09199_),
    .A2(_09384_),
    .B1(_00724_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00727_));
 sky130_fd_sc_hd__o211ai_2 _19536_ (.A1(_09199_),
    .A2(_09384_),
    .B1(_00724_),
    .C1(_00725_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_2 _19537_ (.A(_00726_),
    .B(_00728_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00729_));
 sky130_fd_sc_hd__a31oi_2 _19538_ (.A1(_00631_),
    .A2(_00634_),
    .A3(_00682_),
    .B1(_00680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00731_));
 sky130_fd_sc_hd__a31o_2 _19539_ (.A1(_00631_),
    .A2(_00634_),
    .A3(_00682_),
    .B1(_00680_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00732_));
 sky130_fd_sc_hd__nor2_2 _19540_ (.A(_09220_),
    .B(_09373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00733_));
 sky130_fd_sc_hd__and4_2 _19541_ (.A(\b_l[4] ),
    .B(\b_l[5] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00734_));
 sky130_fd_sc_hd__or3_2 _19542_ (.A(_09220_),
    .B(_09373_),
    .C(_10170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00735_));
 sky130_fd_sc_hd__a22oi_2 _19543_ (.A1(\b_l[5] ),
    .A2(\a_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00736_));
 sky130_fd_sc_hd__nor2_2 _19544_ (.A(_00734_),
    .B(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00737_));
 sky130_fd_sc_hd__a31o_2 _19545_ (.A1(\b_l[4] ),
    .A2(\a_l[14] ),
    .A3(_00733_),
    .B1(_00736_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00738_));
 sky130_fd_sc_hd__a22oi_2 _19546_ (.A1(_10170_),
    .A2(_00637_),
    .B1(_00639_),
    .B2(_00636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00739_));
 sky130_fd_sc_hd__a22o_2 _19547_ (.A1(_10170_),
    .A2(_00637_),
    .B1(_00639_),
    .B2(_00636_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_2 _19548_ (.A(_09264_),
    .B(_09297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00742_));
 sky130_fd_sc_hd__nand2_2 _19549_ (.A(\b_l[8] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_2 _19550_ (.A(\b_l[6] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00744_));
 sky130_fd_sc_hd__and4_2 _19551_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[12] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00745_));
 sky130_fd_sc_hd__nand4_2 _19552_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[12] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00746_));
 sky130_fd_sc_hd__a22oi_2 _19553_ (.A1(\b_l[7] ),
    .A2(\a_l[12] ),
    .B1(\a_l[13] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2_2 _19554_ (.A(_00653_),
    .B(_00744_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00748_));
 sky130_fd_sc_hd__nand2_2 _19555_ (.A(_00746_),
    .B(_00748_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00749_));
 sky130_fd_sc_hd__o2bb2ai_2 _19556_ (.A1_N(_00746_),
    .A2_N(_00748_),
    .B1(_09264_),
    .B2(_09297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00750_));
 sky130_fd_sc_hd__nand4_2 _19557_ (.A(_00748_),
    .B(\a_l[11] ),
    .C(\b_l[8] ),
    .D(_00746_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00751_));
 sky130_fd_sc_hd__a21oi_2 _19558_ (.A1(_00746_),
    .A2(_00748_),
    .B1(_00743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00752_));
 sky130_fd_sc_hd__nand2_2 _19559_ (.A(_00749_),
    .B(_00742_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00753_));
 sky130_fd_sc_hd__o32a_2 _19560_ (.A1(_09319_),
    .A2(_09340_),
    .A3(_04260_),
    .B1(_09297_),
    .B2(_09264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00754_));
 sky130_fd_sc_hd__o21ai_2 _19561_ (.A1(_00653_),
    .A2(_00744_),
    .B1(_00743_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00755_));
 sky130_fd_sc_hd__o21ai_2 _19562_ (.A1(_00747_),
    .A2(_00755_),
    .B1(_00740_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00756_));
 sky130_fd_sc_hd__a21oi_2 _19563_ (.A1(_00750_),
    .A2(_00751_),
    .B1(_00739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00757_));
 sky130_fd_sc_hd__o211ai_2 _19564_ (.A1(_00755_),
    .A2(_00747_),
    .B1(_00740_),
    .C1(_00753_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00758_));
 sky130_fd_sc_hd__o31a_2 _19565_ (.A1(_00747_),
    .A2(_00743_),
    .A3(_00745_),
    .B1(_00739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00759_));
 sky130_fd_sc_hd__nand3_2 _19566_ (.A(_00750_),
    .B(_00751_),
    .C(_00739_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00760_));
 sky130_fd_sc_hd__o21ai_2 _19567_ (.A1(_00752_),
    .A2(_00756_),
    .B1(_00760_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00761_));
 sky130_fd_sc_hd__o32a_2 _19568_ (.A1(_09264_),
    .A2(_09286_),
    .A3(_00651_),
    .B1(_00653_),
    .B2(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00763_));
 sky130_fd_sc_hd__o32ai_2 _19569_ (.A1(_09264_),
    .A2(_09286_),
    .A3(_00651_),
    .B1(_00653_),
    .B2(_00455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00764_));
 sky130_fd_sc_hd__a21oi_2 _19570_ (.A1(_00758_),
    .A2(_00760_),
    .B1(_00764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_2 _19571_ (.A(_00761_),
    .B(_00763_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00766_));
 sky130_fd_sc_hd__o211a_2 _19572_ (.A1(_00752_),
    .A2(_00756_),
    .B1(_00760_),
    .C1(_00764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00767_));
 sky130_fd_sc_hd__o211ai_2 _19573_ (.A1(_00752_),
    .A2(_00756_),
    .B1(_00760_),
    .C1(_00764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2_2 _19574_ (.A(_00766_),
    .B(_00768_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00769_));
 sky130_fd_sc_hd__o22ai_2 _19575_ (.A1(_00734_),
    .A2(_00736_),
    .B1(_00765_),
    .B2(_00767_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00770_));
 sky130_fd_sc_hd__nand3_2 _19576_ (.A(_00766_),
    .B(_00768_),
    .C(_00737_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_2 _19577_ (.A(_00770_),
    .B(_00771_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00772_));
 sky130_fd_sc_hd__a21boi_2 _19578_ (.A1(_00671_),
    .A2(_00673_),
    .B1_N(_00643_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00774_));
 sky130_fd_sc_hd__nand3_2 _19579_ (.A(_00643_),
    .B(_00667_),
    .C(_00669_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_2 _19580_ (.A(_00645_),
    .B(_00775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00776_));
 sky130_fd_sc_hd__o2bb2ai_2 _19581_ (.A1_N(_00770_),
    .A2_N(_00771_),
    .B1(_00774_),
    .B2(_00646_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00777_));
 sky130_fd_sc_hd__nor2_2 _19582_ (.A(_00776_),
    .B(_00772_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00778_));
 sky130_fd_sc_hd__nand4_2 _19583_ (.A(_00645_),
    .B(_00770_),
    .C(_00771_),
    .D(_00775_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_2 _19584_ (.A(_00777_),
    .B(_00779_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00780_));
 sky130_fd_sc_hd__o21ai_2 _19585_ (.A1(_00459_),
    .A2(_00663_),
    .B1(_00661_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_2 _19586_ (.A(_00662_),
    .B(_00781_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00782_));
 sky130_fd_sc_hd__a21boi_2 _19587_ (.A1(_00661_),
    .A2(_00665_),
    .B1_N(_00662_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00783_));
 sky130_fd_sc_hd__nand2_2 _19588_ (.A(\a_l[6] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00785_));
 sky130_fd_sc_hd__nand2_2 _19589_ (.A(\a_l[7] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00786_));
 sky130_fd_sc_hd__and3_2 _19590_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00787_));
 sky130_fd_sc_hd__nand4_2 _19591_ (.A(\a_l[6] ),
    .B(\a_l[7] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00788_));
 sky130_fd_sc_hd__nand2_2 _19592_ (.A(_00785_),
    .B(_00786_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00789_));
 sky130_fd_sc_hd__and4_2 _19593_ (.A(_00789_),
    .B(\b_l[14] ),
    .C(\a_l[5] ),
    .D(_00788_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00790_));
 sky130_fd_sc_hd__or4b_2 _19594_ (.A(_09210_),
    .B(_09362_),
    .C(_00787_),
    .D_N(_00789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00791_));
 sky130_fd_sc_hd__a22oi_2 _19595_ (.A1(\a_l[5] ),
    .A2(\b_l[14] ),
    .B1(_00788_),
    .B2(_00789_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00792_));
 sky130_fd_sc_hd__nor2_2 _19596_ (.A(_00790_),
    .B(_00792_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00793_));
 sky130_fd_sc_hd__a21oi_2 _19597_ (.A1(_00596_),
    .A2(_00597_),
    .B1(_00595_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00794_));
 sky130_fd_sc_hd__a21o_2 _19598_ (.A1(_00595_),
    .A2(_00601_),
    .B1(_00598_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00796_));
 sky130_fd_sc_hd__nand2_2 _19599_ (.A(\a_l[9] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_2 _19600_ (.A(\b_l[9] ),
    .B(\a_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00798_));
 sky130_fd_sc_hd__a22oi_2 _19601_ (.A1(\b_l[9] ),
    .A2(\a_l[10] ),
    .B1(\b_l[10] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_2 _19602_ (.A(_00797_),
    .B(_00798_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00800_));
 sky130_fd_sc_hd__nand4_2 _19603_ (.A(\a_l[9] ),
    .B(\b_l[9] ),
    .C(\a_l[10] ),
    .D(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00801_));
 sky130_fd_sc_hd__nand2_2 _19604_ (.A(\a_l[8] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00802_));
 sky130_fd_sc_hd__nand4_2 _19605_ (.A(_00800_),
    .B(_00801_),
    .C(\a_l[8] ),
    .D(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00803_));
 sky130_fd_sc_hd__o2bb2ai_2 _19606_ (.A1_N(_00800_),
    .A2_N(_00801_),
    .B1(_09253_),
    .B2(_09308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00804_));
 sky130_fd_sc_hd__a21o_2 _19607_ (.A1(_00800_),
    .A2(_00801_),
    .B1(_00802_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00805_));
 sky130_fd_sc_hd__o211ai_2 _19608_ (.A1(_09253_),
    .A2(_09308_),
    .B1(_00800_),
    .C1(_00801_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00807_));
 sky130_fd_sc_hd__o211ai_2 _19609_ (.A1(_00600_),
    .A2(_00794_),
    .B1(_00803_),
    .C1(_00804_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00808_));
 sky130_fd_sc_hd__inv_2 _19610_ (.A(_00808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00809_));
 sky130_fd_sc_hd__and3_2 _19611_ (.A(_00805_),
    .B(_00807_),
    .C(_00796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00810_));
 sky130_fd_sc_hd__nand3_2 _19612_ (.A(_00805_),
    .B(_00807_),
    .C(_00796_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_2 _19613_ (.A(_00808_),
    .B(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_2 _19614_ (.A(_00793_),
    .B(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00813_));
 sky130_fd_sc_hd__o21ai_2 _19615_ (.A1(_00790_),
    .A2(_00792_),
    .B1(_00812_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00814_));
 sky130_fd_sc_hd__o211ai_2 _19616_ (.A1(_00790_),
    .A2(_00792_),
    .B1(_00808_),
    .C1(_00811_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00815_));
 sky130_fd_sc_hd__nand2_2 _19617_ (.A(_00812_),
    .B(_00793_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00816_));
 sky130_fd_sc_hd__nand3_2 _19618_ (.A(_00783_),
    .B(_00815_),
    .C(_00816_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00817_));
 sky130_fd_sc_hd__o211a_2 _19619_ (.A1(_00809_),
    .A2(_00813_),
    .B1(_00782_),
    .C1(_00814_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00818_));
 sky130_fd_sc_hd__o211ai_2 _19620_ (.A1(_00809_),
    .A2(_00813_),
    .B1(_00814_),
    .C1(_00782_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00819_));
 sky130_fd_sc_hd__o21a_2 _19621_ (.A1(_00617_),
    .A2(_00618_),
    .B1(_00607_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00820_));
 sky130_fd_sc_hd__o21ai_2 _19622_ (.A1(_00606_),
    .A2(_00621_),
    .B1(_00608_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00821_));
 sky130_fd_sc_hd__a21oi_2 _19623_ (.A1(_00607_),
    .A2(_00623_),
    .B1(_00609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00822_));
 sky130_fd_sc_hd__o2bb2ai_2 _19624_ (.A1_N(_00817_),
    .A2_N(_00819_),
    .B1(_00820_),
    .B2(_00609_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00823_));
 sky130_fd_sc_hd__a31oi_2 _19625_ (.A1(_00783_),
    .A2(_00815_),
    .A3(_00816_),
    .B1(_00821_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_2 _19626_ (.A(_00817_),
    .B(_00822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00825_));
 sky130_fd_sc_hd__nand3_2 _19627_ (.A(_00817_),
    .B(_00819_),
    .C(_00822_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00826_));
 sky130_fd_sc_hd__o21ai_2 _19628_ (.A1(_00818_),
    .A2(_00825_),
    .B1(_00823_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00828_));
 sky130_fd_sc_hd__a22oi_2 _19629_ (.A1(_00777_),
    .A2(_00779_),
    .B1(_00823_),
    .B2(_00826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00829_));
 sky130_fd_sc_hd__nand2_2 _19630_ (.A(_00780_),
    .B(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00830_));
 sky130_fd_sc_hd__nand3_2 _19631_ (.A(_00777_),
    .B(_00823_),
    .C(_00826_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00831_));
 sky130_fd_sc_hd__o211ai_2 _19632_ (.A1(_00818_),
    .A2(_00825_),
    .B1(_00823_),
    .C1(_00780_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00832_));
 sky130_fd_sc_hd__nand3_2 _19633_ (.A(_00777_),
    .B(_00779_),
    .C(_00828_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00833_));
 sky130_fd_sc_hd__o21ai_2 _19634_ (.A1(_00780_),
    .A2(_00828_),
    .B1(_00732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00834_));
 sky130_fd_sc_hd__o211ai_2 _19635_ (.A1(_00778_),
    .A2(_00831_),
    .B1(_00830_),
    .C1(_00732_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00835_));
 sky130_fd_sc_hd__nand3_2 _19636_ (.A(_00832_),
    .B(_00833_),
    .C(_00731_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00836_));
 sky130_fd_sc_hd__o211ai_2 _19637_ (.A1(_00829_),
    .A2(_00834_),
    .B1(_00836_),
    .C1(_00729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00837_));
 sky130_fd_sc_hd__a21o_2 _19638_ (.A1(_00835_),
    .A2(_00836_),
    .B1(_00729_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00839_));
 sky130_fd_sc_hd__a22o_2 _19639_ (.A1(_00726_),
    .A2(_00728_),
    .B1(_00835_),
    .B2(_00836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00840_));
 sky130_fd_sc_hd__nand4_2 _19640_ (.A(_00726_),
    .B(_00728_),
    .C(_00835_),
    .D(_00836_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_2 _19641_ (.A(_00837_),
    .B(_00839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00842_));
 sky130_fd_sc_hd__nand3_2 _19642_ (.A(_00721_),
    .B(_00837_),
    .C(_00839_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00843_));
 sky130_fd_sc_hd__nand3_2 _19643_ (.A(_00840_),
    .B(_00841_),
    .C(_00720_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00844_));
 sky130_fd_sc_hd__a21bo_2 _19644_ (.A1(_00843_),
    .A2(_00844_),
    .B1_N(_00717_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00845_));
 sky130_fd_sc_hd__o21ai_2 _19645_ (.A1(_00584_),
    .A2(_00587_),
    .B1(_00844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00846_));
 sky130_fd_sc_hd__o211ai_2 _19646_ (.A1(_00584_),
    .A2(_00587_),
    .B1(_00843_),
    .C1(_00844_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00847_));
 sky130_fd_sc_hd__nand2_2 _19647_ (.A(_00845_),
    .B(_00847_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00848_));
 sky130_fd_sc_hd__o21ai_2 _19648_ (.A1(_00549_),
    .A2(_00703_),
    .B1(_00701_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00850_));
 sky130_fd_sc_hd__nand2_2 _19649_ (.A(_00702_),
    .B(_00850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00851_));
 sky130_fd_sc_hd__a22oi_2 _19650_ (.A1(_00845_),
    .A2(_00847_),
    .B1(_00850_),
    .B2(_00702_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00852_));
 sky130_fd_sc_hd__nand2_2 _19651_ (.A(_00848_),
    .B(_00851_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00853_));
 sky130_fd_sc_hd__nand4_2 _19652_ (.A(_00702_),
    .B(_00845_),
    .C(_00847_),
    .D(_00850_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_2 _19653_ (.A(_00853_),
    .B(_00854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_2 _19654_ (.A(_00708_),
    .B(_00716_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00856_));
 sky130_fd_sc_hd__a31o_2 _19655_ (.A1(_00708_),
    .A2(_00716_),
    .A3(_00855_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00857_));
 sky130_fd_sc_hd__a31oi_2 _19656_ (.A1(_00853_),
    .A2(_00854_),
    .A3(_00856_),
    .B1(_00857_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00389_));
 sky130_fd_sc_hd__o21ai_2 _19657_ (.A1(_00720_),
    .A2(_00842_),
    .B1(_00846_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00858_));
 sky130_fd_sc_hd__o2bb2ai_2 _19658_ (.A1_N(_00729_),
    .A2_N(_00836_),
    .B1(_00834_),
    .B2(_00829_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00860_));
 sky130_fd_sc_hd__a21boi_2 _19659_ (.A1(_00729_),
    .A2(_00836_),
    .B1_N(_00835_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00861_));
 sky130_fd_sc_hd__o22a_2 _19660_ (.A1(_00787_),
    .A2(_00790_),
    .B1(_00818_),
    .B2(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00862_));
 sky130_fd_sc_hd__o22ai_2 _19661_ (.A1(_00787_),
    .A2(_00790_),
    .B1(_00818_),
    .B2(_00824_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00863_));
 sky130_fd_sc_hd__o2111ai_2 _19662_ (.A1(_05044_),
    .A2(_06761_),
    .B1(_00791_),
    .C1(_00819_),
    .D1(_00825_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00864_));
 sky130_fd_sc_hd__a22o_2 _19663_ (.A1(\a_l[5] ),
    .A2(\b_l[15] ),
    .B1(_00863_),
    .B2(_00864_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00865_));
 sky130_fd_sc_hd__nand4_2 _19664_ (.A(_00863_),
    .B(_00864_),
    .C(\a_l[5] ),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00866_));
 sky130_fd_sc_hd__nand2_2 _19665_ (.A(_00865_),
    .B(_00866_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00867_));
 sky130_fd_sc_hd__a31oi_2 _19666_ (.A1(_00777_),
    .A2(_00823_),
    .A3(_00826_),
    .B1(_00778_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00868_));
 sky130_fd_sc_hd__o21ai_2 _19667_ (.A1(_00772_),
    .A2(_00776_),
    .B1(_00831_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00869_));
 sky130_fd_sc_hd__nand2_2 _19668_ (.A(\b_l[8] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_2 _19669_ (.A(\b_l[7] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_2 _19670_ (.A(\b_l[7] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_2 _19671_ (.A(\b_l[6] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00874_));
 sky130_fd_sc_hd__nand4_2 _19672_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[13] ),
    .D(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00875_));
 sky130_fd_sc_hd__a22oi_2 _19673_ (.A1(\b_l[7] ),
    .A2(\a_l[13] ),
    .B1(\a_l[14] ),
    .B2(\b_l[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_2 _19674_ (.A(_00873_),
    .B(_00874_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00877_));
 sky130_fd_sc_hd__o2bb2ai_2 _19675_ (.A1_N(_00875_),
    .A2_N(_00877_),
    .B1(_09264_),
    .B2(_09319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00878_));
 sky130_fd_sc_hd__a41o_2 _19676_ (.A1(\b_l[6] ),
    .A2(\b_l[7] ),
    .A3(\a_l[13] ),
    .A4(\a_l[14] ),
    .B1(_00871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00879_));
 sky130_fd_sc_hd__nand4_2 _19677_ (.A(_00877_),
    .B(\a_l[12] ),
    .C(\b_l[8] ),
    .D(_00875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_2 _19678_ (.A(_00878_),
    .B(_00880_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00881_));
 sky130_fd_sc_hd__a21oi_2 _19679_ (.A1(_00878_),
    .A2(_00880_),
    .B1(_00734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_2 _19680_ (.A(_00881_),
    .B(_00735_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00883_));
 sky130_fd_sc_hd__o211a_2 _19681_ (.A1(_00876_),
    .A2(_00879_),
    .B1(_00734_),
    .C1(_00878_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00884_));
 sky130_fd_sc_hd__nand3_2 _19682_ (.A(_00878_),
    .B(_00880_),
    .C(_00734_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00885_));
 sky130_fd_sc_hd__a31o_2 _19683_ (.A1(\b_l[8] ),
    .A2(_00748_),
    .A3(\a_l[11] ),
    .B1(_00745_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00886_));
 sky130_fd_sc_hd__o32a_2 _19684_ (.A1(_09319_),
    .A2(_09340_),
    .A3(_04260_),
    .B1(_00743_),
    .B2(_00747_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00887_));
 sky130_fd_sc_hd__o22ai_2 _19685_ (.A1(_00747_),
    .A2(_00754_),
    .B1(_00882_),
    .B2(_00884_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00888_));
 sky130_fd_sc_hd__nand3_2 _19686_ (.A(_00883_),
    .B(_00885_),
    .C(_00886_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00889_));
 sky130_fd_sc_hd__a21oi_2 _19687_ (.A1(_00881_),
    .A2(_00886_),
    .B1(_00733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00890_));
 sky130_fd_sc_hd__o31ai_2 _19688_ (.A1(_00882_),
    .A2(_00884_),
    .A3(_00886_),
    .B1(_00890_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00892_));
 sky130_fd_sc_hd__nand4_2 _19689_ (.A(_00888_),
    .B(_00889_),
    .C(\b_l[5] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00893_));
 sky130_fd_sc_hd__o2bb2ai_2 _19690_ (.A1_N(_00892_),
    .A2_N(_00893_),
    .B1(_00738_),
    .B2(_00769_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00894_));
 sky130_fd_sc_hd__nand3b_2 _19691_ (.A_N(_00771_),
    .B(_00892_),
    .C(_00893_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00895_));
 sky130_fd_sc_hd__nand2_2 _19692_ (.A(_00894_),
    .B(_00895_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00896_));
 sky130_fd_sc_hd__a22oi_2 _19693_ (.A1(_00759_),
    .A2(_00750_),
    .B1(_00758_),
    .B2(_00764_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00897_));
 sky130_fd_sc_hd__o2bb2ai_2 _19694_ (.A1_N(_00750_),
    .A2_N(_00759_),
    .B1(_00763_),
    .B2(_00757_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2_2 _19695_ (.A(\a_l[7] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_2 _19696_ (.A(\a_l[8] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00900_));
 sky130_fd_sc_hd__and4_2 _19697_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00901_));
 sky130_fd_sc_hd__nand4_2 _19698_ (.A(\a_l[7] ),
    .B(\a_l[8] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00903_));
 sky130_fd_sc_hd__a22oi_2 _19699_ (.A1(\a_l[8] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_2 _19700_ (.A(_00899_),
    .B(_00900_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_2 _19701_ (.A(\a_l[6] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00906_));
 sky130_fd_sc_hd__and4_2 _19702_ (.A(_00905_),
    .B(\b_l[14] ),
    .C(\a_l[6] ),
    .D(_00903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00907_));
 sky130_fd_sc_hd__o22a_2 _19703_ (.A1(_09231_),
    .A2(_09362_),
    .B1(_00901_),
    .B2(_00904_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00908_));
 sky130_fd_sc_hd__and3_2 _19704_ (.A(_00903_),
    .B(_00905_),
    .C(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00909_));
 sky130_fd_sc_hd__a21oi_2 _19705_ (.A1(_00903_),
    .A2(_00905_),
    .B1(_00906_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00910_));
 sky130_fd_sc_hd__and2_2 _19706_ (.A(\a_l[9] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00911_));
 sky130_fd_sc_hd__nand2_2 _19707_ (.A(\a_l[9] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_2 _19708_ (.A(\a_l[10] ),
    .B(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_2 _19709_ (.A(\b_l[9] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_2 _19710_ (.A(\b_l[9] ),
    .B(\a_l[10] ),
    .C(\b_l[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00916_));
 sky130_fd_sc_hd__nand4_2 _19711_ (.A(\b_l[9] ),
    .B(\a_l[10] ),
    .C(\b_l[10] ),
    .D(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00917_));
 sky130_fd_sc_hd__a22oi_2 _19712_ (.A1(\a_l[10] ),
    .A2(\b_l[10] ),
    .B1(\a_l[11] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00918_));
 sky130_fd_sc_hd__nand2_2 _19713_ (.A(_00914_),
    .B(_00915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00919_));
 sky130_fd_sc_hd__o21ai_2 _19714_ (.A1(_09297_),
    .A2(_00916_),
    .B1(_00919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00920_));
 sky130_fd_sc_hd__o21ai_2 _19715_ (.A1(_09275_),
    .A2(_09308_),
    .B1(_00920_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00921_));
 sky130_fd_sc_hd__a41o_2 _19716_ (.A1(\b_l[9] ),
    .A2(\a_l[10] ),
    .A3(\b_l[10] ),
    .A4(\a_l[11] ),
    .B1(_00912_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00922_));
 sky130_fd_sc_hd__a21o_2 _19717_ (.A1(_00801_),
    .A2(_00802_),
    .B1(_00799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00923_));
 sky130_fd_sc_hd__a21oi_2 _19718_ (.A1(_00801_),
    .A2(_00802_),
    .B1(_00799_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00925_));
 sky130_fd_sc_hd__o211a_2 _19719_ (.A1(_00918_),
    .A2(_00922_),
    .B1(_00925_),
    .C1(_00921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00926_));
 sky130_fd_sc_hd__o211ai_2 _19720_ (.A1(_00918_),
    .A2(_00922_),
    .B1(_00925_),
    .C1(_00921_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00927_));
 sky130_fd_sc_hd__o221ai_2 _19721_ (.A1(_09275_),
    .A2(_09308_),
    .B1(_00916_),
    .B2(_09297_),
    .C1(_00919_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_2 _19722_ (.A(_00920_),
    .B(_00911_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00929_));
 sky130_fd_sc_hd__and3_2 _19723_ (.A(_00929_),
    .B(_00923_),
    .C(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00930_));
 sky130_fd_sc_hd__nand3_2 _19724_ (.A(_00929_),
    .B(_00923_),
    .C(_00928_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_2 _19725_ (.A(_00927_),
    .B(_00931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00932_));
 sky130_fd_sc_hd__o211ai_2 _19726_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00927_),
    .C1(_00931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00933_));
 sky130_fd_sc_hd__o21ai_2 _19727_ (.A1(_00909_),
    .A2(_00910_),
    .B1(_00932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00934_));
 sky130_fd_sc_hd__o21ai_2 _19728_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00932_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00936_));
 sky130_fd_sc_hd__o21ai_2 _19729_ (.A1(_00909_),
    .A2(_00910_),
    .B1(_00931_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00937_));
 sky130_fd_sc_hd__o211a_2 _19730_ (.A1(_00937_),
    .A2(_00926_),
    .B1(_00898_),
    .C1(_00936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00938_));
 sky130_fd_sc_hd__o211ai_2 _19731_ (.A1(_00937_),
    .A2(_00926_),
    .B1(_00898_),
    .C1(_00936_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00939_));
 sky130_fd_sc_hd__nand3_2 _19732_ (.A(_00934_),
    .B(_00897_),
    .C(_00933_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00940_));
 sky130_fd_sc_hd__o21a_2 _19733_ (.A1(_00790_),
    .A2(_00792_),
    .B1(_00808_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00941_));
 sky130_fd_sc_hd__a21o_2 _19734_ (.A1(_00793_),
    .A2(_00811_),
    .B1(_00809_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00942_));
 sky130_fd_sc_hd__nand2_2 _19735_ (.A(_00940_),
    .B(_00942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00943_));
 sky130_fd_sc_hd__nand3_2 _19736_ (.A(_00939_),
    .B(_00940_),
    .C(_00942_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00944_));
 sky130_fd_sc_hd__o2bb2ai_2 _19737_ (.A1_N(_00939_),
    .A2_N(_00940_),
    .B1(_00941_),
    .B2(_00810_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00945_));
 sky130_fd_sc_hd__o21ai_2 _19738_ (.A1(_00810_),
    .A2(_00941_),
    .B1(_00939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00946_));
 sky130_fd_sc_hd__o211ai_2 _19739_ (.A1(_00810_),
    .A2(_00941_),
    .B1(_00940_),
    .C1(_00939_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00947_));
 sky130_fd_sc_hd__a22o_2 _19740_ (.A1(_00808_),
    .A2(_00813_),
    .B1(_00939_),
    .B2(_00940_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00948_));
 sky130_fd_sc_hd__nand4_2 _19741_ (.A(_00894_),
    .B(_00895_),
    .C(_00944_),
    .D(_00945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00949_));
 sky130_fd_sc_hd__nand3_2 _19742_ (.A(_00896_),
    .B(_00947_),
    .C(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00950_));
 sky130_fd_sc_hd__nand4_2 _19743_ (.A(_00894_),
    .B(_00895_),
    .C(_00947_),
    .D(_00948_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00951_));
 sky130_fd_sc_hd__nand3_2 _19744_ (.A(_00896_),
    .B(_00944_),
    .C(_00945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00952_));
 sky130_fd_sc_hd__nand3_2 _19745_ (.A(_00869_),
    .B(_00949_),
    .C(_00950_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00953_));
 sky130_fd_sc_hd__a21oi_2 _19746_ (.A1(_00949_),
    .A2(_00950_),
    .B1(_00869_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_2 _19747_ (.A(_00868_),
    .B(_00951_),
    .C(_00952_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00955_));
 sky130_fd_sc_hd__a21o_2 _19748_ (.A1(_00953_),
    .A2(_00955_),
    .B1(_00867_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00957_));
 sky130_fd_sc_hd__nand3_2 _19749_ (.A(_00867_),
    .B(_00953_),
    .C(_00955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00958_));
 sky130_fd_sc_hd__nand4_2 _19750_ (.A(_00865_),
    .B(_00866_),
    .C(_00953_),
    .D(_00955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00959_));
 sky130_fd_sc_hd__a22o_2 _19751_ (.A1(_00865_),
    .A2(_00866_),
    .B1(_00953_),
    .B2(_00955_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00960_));
 sky130_fd_sc_hd__nand3_2 _19752_ (.A(_00861_),
    .B(_00957_),
    .C(_00958_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00961_));
 sky130_fd_sc_hd__a21oi_2 _19753_ (.A1(_00957_),
    .A2(_00958_),
    .B1(_00861_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00962_));
 sky130_fd_sc_hd__nand3_2 _19754_ (.A(_00960_),
    .B(_00860_),
    .C(_00959_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00963_));
 sky130_fd_sc_hd__and2_2 _19755_ (.A(_00725_),
    .B(_00727_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00964_));
 sky130_fd_sc_hd__a22o_2 _19756_ (.A1(_00725_),
    .A2(_00727_),
    .B1(_00961_),
    .B2(_00963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00965_));
 sky130_fd_sc_hd__nand4_2 _19757_ (.A(_00725_),
    .B(_00727_),
    .C(_00961_),
    .D(_00963_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00966_));
 sky130_fd_sc_hd__a21o_2 _19758_ (.A1(_00965_),
    .A2(_00966_),
    .B1(_00858_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00968_));
 sky130_fd_sc_hd__nand3_2 _19759_ (.A(_00858_),
    .B(_00965_),
    .C(_00966_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_2 _19760_ (.A(_00968_),
    .B(_00969_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00970_));
 sky130_fd_sc_hd__o21ai_2 _19761_ (.A1(_00708_),
    .A2(_00852_),
    .B1(_00854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00971_));
 sky130_fd_sc_hd__nor2_2 _19762_ (.A(_00710_),
    .B(_00855_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00972_));
 sky130_fd_sc_hd__nand4_2 _19763_ (.A(_00707_),
    .B(_00708_),
    .C(_00853_),
    .D(_00854_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00973_));
 sky130_fd_sc_hd__nor2_2 _19764_ (.A(_00712_),
    .B(_00973_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_2 _19765_ (.A(_10004_),
    .B(_00974_),
    .C(_10002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00975_));
 sky130_fd_sc_hd__a21oi_2 _19766_ (.A1(_00972_),
    .A2(_00713_),
    .B1(_00971_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00976_));
 sky130_fd_sc_hd__o311a_2 _19767_ (.A1(_10005_),
    .A2(_00712_),
    .A3(_00973_),
    .B1(_00976_),
    .C1(_00970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00977_));
 sky130_fd_sc_hd__a21oi_2 _19768_ (.A1(_00975_),
    .A2(_00976_),
    .B1(_00970_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00979_));
 sky130_fd_sc_hd__nor3_2 _19769_ (.A(rst),
    .B(_00977_),
    .C(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00390_));
 sky130_fd_sc_hd__a21oi_2 _19770_ (.A1(_00867_),
    .A2(_00953_),
    .B1(_00954_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00980_));
 sky130_fd_sc_hd__and2_2 _19771_ (.A(\b_l[8] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00981_));
 sky130_fd_sc_hd__nand2_2 _19772_ (.A(\b_l[6] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_2 _19773_ (.A(_00872_),
    .B(_00982_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00983_));
 sky130_fd_sc_hd__nand4_2 _19774_ (.A(\b_l[6] ),
    .B(\b_l[7] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00984_));
 sky130_fd_sc_hd__o2bb2a_2 _19775_ (.A1_N(_00983_),
    .A2_N(_00984_),
    .B1(_09264_),
    .B2(_09340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00985_));
 sky130_fd_sc_hd__o2bb2ai_2 _19776_ (.A1_N(_00983_),
    .A2_N(_00984_),
    .B1(_09264_),
    .B2(_09340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00986_));
 sky130_fd_sc_hd__nand3_2 _19777_ (.A(_00983_),
    .B(_00984_),
    .C(_00981_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00987_));
 sky130_fd_sc_hd__o21ai_2 _19778_ (.A1(_00744_),
    .A2(_00872_),
    .B1(_00871_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00989_));
 sky130_fd_sc_hd__o21ai_2 _19779_ (.A1(_00871_),
    .A2(_00876_),
    .B1(_00875_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00990_));
 sky130_fd_sc_hd__a21oi_2 _19780_ (.A1(_00986_),
    .A2(_00987_),
    .B1(_00990_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00991_));
 sky130_fd_sc_hd__and3_2 _19781_ (.A(_00877_),
    .B(_00987_),
    .C(_00989_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00992_));
 sky130_fd_sc_hd__nand2_2 _19782_ (.A(_00990_),
    .B(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00993_));
 sky130_fd_sc_hd__and3_2 _19783_ (.A(_00986_),
    .B(_00990_),
    .C(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00994_));
 sky130_fd_sc_hd__a21oi_2 _19784_ (.A1(_00992_),
    .A2(_00986_),
    .B1(_00991_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00995_));
 sky130_fd_sc_hd__and4_2 _19785_ (.A(_00888_),
    .B(_00995_),
    .C(_00889_),
    .D(_00733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00996_));
 sky130_fd_sc_hd__nand4_2 _19786_ (.A(_00888_),
    .B(_00995_),
    .C(_00889_),
    .D(_00733_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00997_));
 sky130_fd_sc_hd__a31oi_2 _19787_ (.A1(_00888_),
    .A2(_00889_),
    .A3(_00733_),
    .B1(_00995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00998_));
 sky130_fd_sc_hd__a31o_2 _19788_ (.A1(_00888_),
    .A2(_00889_),
    .A3(_00733_),
    .B1(_00995_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01000_));
 sky130_fd_sc_hd__nor2_2 _19789_ (.A(_00996_),
    .B(_00998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_2 _19790_ (.A(_00885_),
    .B(_00887_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01002_));
 sky130_fd_sc_hd__o21ai_2 _19791_ (.A1(_00887_),
    .A2(_00882_),
    .B1(_00885_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_2 _19792_ (.A(_00883_),
    .B(_01002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01004_));
 sky130_fd_sc_hd__nand2_2 _19793_ (.A(\a_l[8] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_2 _19794_ (.A(\a_l[9] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01006_));
 sky130_fd_sc_hd__nand4_2 _19795_ (.A(\a_l[8] ),
    .B(\a_l[9] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_2 _19796_ (.A(_01005_),
    .B(_01006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01008_));
 sky130_fd_sc_hd__and4_2 _19797_ (.A(_01008_),
    .B(\b_l[14] ),
    .C(\a_l[7] ),
    .D(_01007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01009_));
 sky130_fd_sc_hd__a22oi_2 _19798_ (.A1(\a_l[7] ),
    .A2(\b_l[14] ),
    .B1(_01007_),
    .B2(_01008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01011_));
 sky130_fd_sc_hd__nor2_2 _19799_ (.A(_01009_),
    .B(_01011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01012_));
 sky130_fd_sc_hd__o21ai_2 _19800_ (.A1(_00912_),
    .A2(_00918_),
    .B1(_00917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01013_));
 sky130_fd_sc_hd__a21boi_2 _19801_ (.A1(_00919_),
    .A2(_00911_),
    .B1_N(_00917_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01014_));
 sky130_fd_sc_hd__and2_2 _19802_ (.A(\a_l[10] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01015_));
 sky130_fd_sc_hd__nand2_2 _19803_ (.A(\a_l[10] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_2 _19804_ (.A(\b_l[10] ),
    .B(\a_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_2 _19805_ (.A(\b_l[9] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01018_));
 sky130_fd_sc_hd__a22o_2 _19806_ (.A1(\b_l[10] ),
    .A2(\a_l[11] ),
    .B1(\a_l[12] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01019_));
 sky130_fd_sc_hd__nand2_2 _19807_ (.A(\b_l[10] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01020_));
 sky130_fd_sc_hd__nand4_2 _19808_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_l[11] ),
    .D(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01022_));
 sky130_fd_sc_hd__o2bb2ai_2 _19809_ (.A1_N(_01017_),
    .A2_N(_01018_),
    .B1(_01020_),
    .B2(_00915_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01023_));
 sky130_fd_sc_hd__o211ai_2 _19810_ (.A1(_00915_),
    .A2(_01020_),
    .B1(_01015_),
    .C1(_01019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01024_));
 sky130_fd_sc_hd__o21ai_2 _19811_ (.A1(_09286_),
    .A2(_09308_),
    .B1(_01023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01025_));
 sky130_fd_sc_hd__nand2_2 _19812_ (.A(_01023_),
    .B(_01015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01026_));
 sky130_fd_sc_hd__o221ai_2 _19813_ (.A1(_09286_),
    .A2(_09308_),
    .B1(_00915_),
    .B2(_01020_),
    .C1(_01019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01027_));
 sky130_fd_sc_hd__nand3_2 _19814_ (.A(_01025_),
    .B(_01013_),
    .C(_01024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01028_));
 sky130_fd_sc_hd__a21oi_2 _19815_ (.A1(_01024_),
    .A2(_01025_),
    .B1(_01013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01029_));
 sky130_fd_sc_hd__nand3_2 _19816_ (.A(_01014_),
    .B(_01026_),
    .C(_01027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_2 _19817_ (.A(_01028_),
    .B(_01030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_2 _19818_ (.A(_01031_),
    .B(_01012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01032_));
 sky130_fd_sc_hd__o21ai_2 _19819_ (.A1(_01009_),
    .A2(_01011_),
    .B1(_01028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01033_));
 sky130_fd_sc_hd__nand3_2 _19820_ (.A(_01012_),
    .B(_01028_),
    .C(_01030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01034_));
 sky130_fd_sc_hd__o21ai_2 _19821_ (.A1(_01009_),
    .A2(_01011_),
    .B1(_01031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01035_));
 sky130_fd_sc_hd__nand3_2 _19822_ (.A(_01035_),
    .B(_01003_),
    .C(_01034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01036_));
 sky130_fd_sc_hd__o211ai_2 _19823_ (.A1(_01033_),
    .A2(_01029_),
    .B1(_01004_),
    .C1(_01032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01037_));
 sky130_fd_sc_hd__o21a_2 _19824_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00927_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01038_));
 sky130_fd_sc_hd__nand2_2 _19825_ (.A(_00927_),
    .B(_00937_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01039_));
 sky130_fd_sc_hd__a22oi_2 _19826_ (.A1(_00927_),
    .A2(_00937_),
    .B1(_01036_),
    .B2(_01037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01040_));
 sky130_fd_sc_hd__a22o_2 _19827_ (.A1(_00927_),
    .A2(_00937_),
    .B1(_01036_),
    .B2(_01037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01041_));
 sky130_fd_sc_hd__nand3b_2 _19828_ (.A_N(_01039_),
    .B(_01037_),
    .C(_01036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01043_));
 sky130_fd_sc_hd__nand3_2 _19829_ (.A(_01036_),
    .B(_01037_),
    .C(_01039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01044_));
 sky130_fd_sc_hd__o2bb2ai_2 _19830_ (.A1_N(_01036_),
    .A2_N(_01037_),
    .B1(_01038_),
    .B2(_00930_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01045_));
 sky130_fd_sc_hd__o211ai_2 _19831_ (.A1(_00996_),
    .A2(_00998_),
    .B1(_01044_),
    .C1(_01045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01046_));
 sky130_fd_sc_hd__nand3_2 _19832_ (.A(_00997_),
    .B(_01041_),
    .C(_01043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01047_));
 sky130_fd_sc_hd__nand3_2 _19833_ (.A(_00997_),
    .B(_01000_),
    .C(_01043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01048_));
 sky130_fd_sc_hd__nand3_2 _19834_ (.A(_01001_),
    .B(_01041_),
    .C(_01043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01049_));
 sky130_fd_sc_hd__o21ai_2 _19835_ (.A1(_01040_),
    .A2(_01048_),
    .B1(_01046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01050_));
 sky130_fd_sc_hd__o211ai_2 _19836_ (.A1(_00943_),
    .A2(_00938_),
    .B1(_00894_),
    .C1(_00945_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01051_));
 sky130_fd_sc_hd__nand2_2 _19837_ (.A(_00895_),
    .B(_01051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_2 _19838_ (.A(_01052_),
    .B(_01050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01054_));
 sky130_fd_sc_hd__nor2_2 _19839_ (.A(_01050_),
    .B(_01052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01055_));
 sky130_fd_sc_hd__nand4_2 _19840_ (.A(_00895_),
    .B(_01046_),
    .C(_01049_),
    .D(_01051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01056_));
 sky130_fd_sc_hd__nand2_2 _19841_ (.A(_01054_),
    .B(_01056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01057_));
 sky130_fd_sc_hd__o31a_2 _19842_ (.A1(_09231_),
    .A2(_09362_),
    .A3(_00904_),
    .B1(_00903_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01058_));
 sky130_fd_sc_hd__nand3_2 _19843_ (.A(_00939_),
    .B(_00943_),
    .C(_01058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01059_));
 sky130_fd_sc_hd__o211ai_2 _19844_ (.A1(_00901_),
    .A2(_00907_),
    .B1(_00940_),
    .C1(_00946_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01060_));
 sky130_fd_sc_hd__o2bb2ai_2 _19845_ (.A1_N(_01059_),
    .A2_N(_01060_),
    .B1(_09231_),
    .B2(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01061_));
 sky130_fd_sc_hd__nand4_2 _19846_ (.A(_01060_),
    .B(\a_l[6] ),
    .C(_01059_),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01062_));
 sky130_fd_sc_hd__and2_2 _19847_ (.A(_01061_),
    .B(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01063_));
 sky130_fd_sc_hd__nand2_2 _19848_ (.A(_01061_),
    .B(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_2 _19849_ (.A(_01054_),
    .B(_01056_),
    .C(_01065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_2 _19850_ (.A(_01057_),
    .B(_01063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01067_));
 sky130_fd_sc_hd__o2111ai_2 _19851_ (.A1(_00954_),
    .A2(_00867_),
    .B1(_00953_),
    .C1(_01066_),
    .D1(_01067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01068_));
 sky130_fd_sc_hd__nand4_2 _19852_ (.A(_01054_),
    .B(_01056_),
    .C(_01061_),
    .D(_01062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_2 _19853_ (.A(_01057_),
    .B(_01065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01070_));
 sky130_fd_sc_hd__nand3_2 _19854_ (.A(_00980_),
    .B(_01069_),
    .C(_01070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_2 _19855_ (.A(_01068_),
    .B(_01071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01072_));
 sky130_fd_sc_hd__a31o_2 _19856_ (.A1(\a_l[5] ),
    .A2(\b_l[15] ),
    .A3(_00864_),
    .B1(_00862_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01073_));
 sky130_fd_sc_hd__inv_2 _19857_ (.A(_01073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01074_));
 sky130_fd_sc_hd__nand2_2 _19858_ (.A(_01072_),
    .B(_01074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01075_));
 sky130_fd_sc_hd__nand3_2 _19859_ (.A(_01068_),
    .B(_01071_),
    .C(_01073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01076_));
 sky130_fd_sc_hd__a21o_2 _19860_ (.A1(_00961_),
    .A2(_00964_),
    .B1(_00962_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01077_));
 sky130_fd_sc_hd__a21oi_2 _19861_ (.A1(_01075_),
    .A2(_01076_),
    .B1(_01077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01078_));
 sky130_fd_sc_hd__a21o_2 _19862_ (.A1(_01075_),
    .A2(_01076_),
    .B1(_01077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01079_));
 sky130_fd_sc_hd__nand3_2 _19863_ (.A(_01077_),
    .B(_01076_),
    .C(_01075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_2 _19864_ (.A(_01079_),
    .B(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01081_));
 sky130_fd_sc_hd__a31oi_2 _19865_ (.A1(_00858_),
    .A2(_00965_),
    .A3(_00966_),
    .B1(_00979_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01082_));
 sky130_fd_sc_hd__o21ai_2 _19866_ (.A1(_01081_),
    .A2(_01082_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_2 _19867_ (.A1(_01081_),
    .A2(_01082_),
    .B1(_01083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00391_));
 sky130_fd_sc_hd__a21boi_2 _19868_ (.A1(_01068_),
    .A2(_01073_),
    .B1_N(_01071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01085_));
 sky130_fd_sc_hd__o21ai_2 _19869_ (.A1(_01065_),
    .A2(_01055_),
    .B1(_01054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01086_));
 sky130_fd_sc_hd__o21a_2 _19870_ (.A1(_01065_),
    .A2(_01055_),
    .B1(_01054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01087_));
 sky130_fd_sc_hd__a31o_2 _19871_ (.A1(\b_l[12] ),
    .A2(\b_l[13] ),
    .A3(_06984_),
    .B1(_01009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01088_));
 sky130_fd_sc_hd__a31o_2 _19872_ (.A1(_01035_),
    .A2(_01003_),
    .A3(_01034_),
    .B1(_01039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01089_));
 sky130_fd_sc_hd__nand3_2 _19873_ (.A(_01037_),
    .B(_01088_),
    .C(_01089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01090_));
 sky130_fd_sc_hd__a21oi_2 _19874_ (.A1(_01037_),
    .A2(_01039_),
    .B1(_01088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01091_));
 sky130_fd_sc_hd__a21oi_2 _19875_ (.A1(_01037_),
    .A2(_01089_),
    .B1(_01088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_2 _19876_ (.A(_01091_),
    .B(_01036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01093_));
 sky130_fd_sc_hd__a22o_2 _19877_ (.A1(\a_l[7] ),
    .A2(\b_l[15] ),
    .B1(_01090_),
    .B2(_01093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01094_));
 sky130_fd_sc_hd__nand4_2 _19878_ (.A(_01093_),
    .B(\a_l[7] ),
    .C(_01090_),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_2 _19879_ (.A(_01094_),
    .B(_01096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01097_));
 sky130_fd_sc_hd__o21a_2 _19880_ (.A1(_00872_),
    .A2(_00982_),
    .B1(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01098_));
 sky130_fd_sc_hd__o21ai_2 _19881_ (.A1(_00872_),
    .A2(_00982_),
    .B1(_00987_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_2 _19882_ (.A(\b_l[8] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01100_));
 sky130_fd_sc_hd__and4_2 _19883_ (.A(\b_l[7] ),
    .B(\b_l[8] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01101_));
 sky130_fd_sc_hd__a22oi_2 _19884_ (.A1(\b_l[8] ),
    .A2(\a_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_2 _19885_ (.A(_01101_),
    .B(_01102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01103_));
 sky130_fd_sc_hd__or2_2 _19886_ (.A(_01101_),
    .B(_01102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01104_));
 sky130_fd_sc_hd__a211o_2 _19887_ (.A1(_00984_),
    .A2(_00987_),
    .B1(_01101_),
    .C1(_01102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01105_));
 sky130_fd_sc_hd__o21ai_2 _19888_ (.A1(_01101_),
    .A2(_01102_),
    .B1(_01098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_2 _19889_ (.A(_01105_),
    .B(_01107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01108_));
 sky130_fd_sc_hd__nand2_2 _19890_ (.A(\a_l[11] ),
    .B(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_2 _19891_ (.A(\b_l[9] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01110_));
 sky130_fd_sc_hd__nand3_2 _19892_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01111_));
 sky130_fd_sc_hd__nand4_2 _19893_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_l[12] ),
    .D(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01112_));
 sky130_fd_sc_hd__a22oi_2 _19894_ (.A1(\b_l[10] ),
    .A2(\a_l[12] ),
    .B1(\a_l[13] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_2 _19895_ (.A(_01020_),
    .B(_01110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01114_));
 sky130_fd_sc_hd__a21bo_2 _19896_ (.A1(_01112_),
    .A2(_01114_),
    .B1_N(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01115_));
 sky130_fd_sc_hd__a41o_2 _19897_ (.A1(\b_l[9] ),
    .A2(\b_l[10] ),
    .A3(\a_l[12] ),
    .A4(\a_l[13] ),
    .B1(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01116_));
 sky130_fd_sc_hd__a22o_2 _19898_ (.A1(_01017_),
    .A2(_01018_),
    .B1(_01022_),
    .B2(_01016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01118_));
 sky130_fd_sc_hd__a22oi_2 _19899_ (.A1(_01017_),
    .A2(_01018_),
    .B1(_01022_),
    .B2(_01016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01119_));
 sky130_fd_sc_hd__o211ai_2 _19900_ (.A1(_01113_),
    .A2(_01116_),
    .B1(_01119_),
    .C1(_01115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01120_));
 sky130_fd_sc_hd__inv_2 _19901_ (.A(_01120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01121_));
 sky130_fd_sc_hd__nand2_2 _19902_ (.A(_01109_),
    .B(_01112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01122_));
 sky130_fd_sc_hd__a21o_2 _19903_ (.A1(_01112_),
    .A2(_01114_),
    .B1(_01109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01123_));
 sky130_fd_sc_hd__o211ai_2 _19904_ (.A1(_01113_),
    .A2(_01122_),
    .B1(_01118_),
    .C1(_01123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_2 _19905_ (.A(\a_l[8] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01125_));
 sky130_fd_sc_hd__a22o_2 _19906_ (.A1(\a_l[10] ),
    .A2(\b_l[12] ),
    .B1(\b_l[13] ),
    .B2(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01126_));
 sky130_fd_sc_hd__and3_2 _19907_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(_05043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01127_));
 sky130_fd_sc_hd__nand4_2 _19908_ (.A(\a_l[9] ),
    .B(\a_l[10] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01129_));
 sky130_fd_sc_hd__a22oi_2 _19909_ (.A1(\a_l[8] ),
    .A2(\b_l[14] ),
    .B1(_01126_),
    .B2(_01129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01130_));
 sky130_fd_sc_hd__and4_2 _19910_ (.A(_01126_),
    .B(_01129_),
    .C(\a_l[8] ),
    .D(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01131_));
 sky130_fd_sc_hd__o311a_2 _19911_ (.A1(_09275_),
    .A2(_09286_),
    .A3(_05044_),
    .B1(_01125_),
    .C1(_01126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01132_));
 sky130_fd_sc_hd__a21oi_2 _19912_ (.A1(_01126_),
    .A2(_01129_),
    .B1(_01125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_2 _19913_ (.A(_01130_),
    .B(_01131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01134_));
 sky130_fd_sc_hd__o2bb2ai_2 _19914_ (.A1_N(_01120_),
    .A2_N(_01124_),
    .B1(_01130_),
    .B2(_01131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01135_));
 sky130_fd_sc_hd__o21ai_2 _19915_ (.A1(_01132_),
    .A2(_01133_),
    .B1(_01124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01136_));
 sky130_fd_sc_hd__inv_2 _19916_ (.A(_01136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01137_));
 sky130_fd_sc_hd__nand3_2 _19917_ (.A(_01134_),
    .B(_01124_),
    .C(_01120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01138_));
 sky130_fd_sc_hd__o2bb2ai_2 _19918_ (.A1_N(_01120_),
    .A2_N(_01124_),
    .B1(_01132_),
    .B2(_01133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01140_));
 sky130_fd_sc_hd__o211ai_2 _19919_ (.A1(_01130_),
    .A2(_01131_),
    .B1(_01120_),
    .C1(_01124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01141_));
 sky130_fd_sc_hd__o211ai_2 _19920_ (.A1(_00993_),
    .A2(_00985_),
    .B1(_01141_),
    .C1(_01140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01142_));
 sky130_fd_sc_hd__nand3_2 _19921_ (.A(_01135_),
    .B(_01138_),
    .C(_00994_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01143_));
 sky130_fd_sc_hd__o31ai_2 _19922_ (.A1(_01009_),
    .A2(_01011_),
    .A3(_01029_),
    .B1(_01028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01144_));
 sky130_fd_sc_hd__o31a_2 _19923_ (.A1(_01009_),
    .A2(_01011_),
    .A3(_01029_),
    .B1(_01028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01145_));
 sky130_fd_sc_hd__a21o_2 _19924_ (.A1(_01142_),
    .A2(_01143_),
    .B1(_01145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01146_));
 sky130_fd_sc_hd__nand3_2 _19925_ (.A(_01142_),
    .B(_01143_),
    .C(_01145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01147_));
 sky130_fd_sc_hd__a21o_2 _19926_ (.A1(_01142_),
    .A2(_01143_),
    .B1(_01144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_2 _19927_ (.A(_01142_),
    .B(_01144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01149_));
 sky130_fd_sc_hd__nand4_2 _19928_ (.A(_01030_),
    .B(_01033_),
    .C(_01142_),
    .D(_01143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01151_));
 sky130_fd_sc_hd__a21oi_2 _19929_ (.A1(_01146_),
    .A2(_01147_),
    .B1(_01108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01152_));
 sky130_fd_sc_hd__nand3b_2 _19930_ (.A_N(_01108_),
    .B(_01148_),
    .C(_01151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01153_));
 sky130_fd_sc_hd__nand3_2 _19931_ (.A(_01108_),
    .B(_01146_),
    .C(_01147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_2 _19932_ (.A(_01153_),
    .B(_01154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01155_));
 sky130_fd_sc_hd__a31o_2 _19933_ (.A1(_00997_),
    .A2(_01041_),
    .A3(_01043_),
    .B1(_00998_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01156_));
 sky130_fd_sc_hd__nand4_2 _19934_ (.A(_01000_),
    .B(_01047_),
    .C(_01153_),
    .D(_01154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_2 _19935_ (.A(_01156_),
    .B(_01155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01158_));
 sky130_fd_sc_hd__inv_2 _19936_ (.A(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01159_));
 sky130_fd_sc_hd__a22o_2 _19937_ (.A1(_01094_),
    .A2(_01096_),
    .B1(_01157_),
    .B2(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01160_));
 sky130_fd_sc_hd__nand4_2 _19938_ (.A(_01094_),
    .B(_01096_),
    .C(_01157_),
    .D(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01162_));
 sky130_fd_sc_hd__nand3_2 _19939_ (.A(_01097_),
    .B(_01157_),
    .C(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01163_));
 sky130_fd_sc_hd__a21o_2 _19940_ (.A1(_01157_),
    .A2(_01158_),
    .B1(_01097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01164_));
 sky130_fd_sc_hd__nand2_2 _19941_ (.A(_01163_),
    .B(_01164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01165_));
 sky130_fd_sc_hd__nand3_2 _19942_ (.A(_01087_),
    .B(_01163_),
    .C(_01164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01166_));
 sky130_fd_sc_hd__inv_2 _19943_ (.A(_01166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01167_));
 sky130_fd_sc_hd__nand3_2 _19944_ (.A(_01160_),
    .B(_01162_),
    .C(_01086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01168_));
 sky130_fd_sc_hd__o21ai_2 _19945_ (.A1(_09231_),
    .A2(_09384_),
    .B1(_01060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_2 _19946_ (.A(_01059_),
    .B(_01169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01170_));
 sky130_fd_sc_hd__inv_2 _19947_ (.A(_01170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01171_));
 sky130_fd_sc_hd__a21o_2 _19948_ (.A1(_01166_),
    .A2(_01168_),
    .B1(_01170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01173_));
 sky130_fd_sc_hd__a31oi_2 _19949_ (.A1(_01160_),
    .A2(_01162_),
    .A3(_01086_),
    .B1(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01174_));
 sky130_fd_sc_hd__a31o_2 _19950_ (.A1(_01160_),
    .A2(_01162_),
    .A3(_01086_),
    .B1(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01175_));
 sky130_fd_sc_hd__and3_2 _19951_ (.A(_01166_),
    .B(_01168_),
    .C(_01170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01176_));
 sky130_fd_sc_hd__nand4_2 _19952_ (.A(_01059_),
    .B(_01166_),
    .C(_01168_),
    .D(_01169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01177_));
 sky130_fd_sc_hd__a21o_2 _19953_ (.A1(_01166_),
    .A2(_01168_),
    .B1(_01171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01178_));
 sky130_fd_sc_hd__nand3b_2 _19954_ (.A_N(_01085_),
    .B(_01177_),
    .C(_01178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_2 _19955_ (.A(_01085_),
    .B(_01173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01180_));
 sky130_fd_sc_hd__o211ai_2 _19956_ (.A1(_01175_),
    .A2(_01167_),
    .B1(_01085_),
    .C1(_01173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01181_));
 sky130_fd_sc_hd__o21a_2 _19957_ (.A1(_01176_),
    .A2(_01180_),
    .B1(_01179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01182_));
 sky130_fd_sc_hd__o21ai_2 _19958_ (.A1(_00969_),
    .A2(_01078_),
    .B1(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01183_));
 sky130_fd_sc_hd__nand4_2 _19959_ (.A(_00968_),
    .B(_00969_),
    .C(_01079_),
    .D(_01080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01184_));
 sky130_fd_sc_hd__a21oi_2 _19960_ (.A1(_00975_),
    .A2(_00976_),
    .B1(_01184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01185_));
 sky130_fd_sc_hd__a211oi_2 _19961_ (.A1(_01179_),
    .A2(_01181_),
    .B1(_01183_),
    .C1(_01185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01186_));
 sky130_fd_sc_hd__o21ai_2 _19962_ (.A1(_01183_),
    .A2(_01185_),
    .B1(_01182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01187_));
 sky130_fd_sc_hd__nor3b_2 _19963_ (.A(rst),
    .B(_01186_),
    .C_N(_01187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00392_));
 sky130_fd_sc_hd__a21boi_2 _19964_ (.A1(_01094_),
    .A2(_01096_),
    .B1_N(_01157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01188_));
 sky130_fd_sc_hd__a21boi_2 _19965_ (.A1(_01097_),
    .A2(_01157_),
    .B1_N(_01158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_2 _19966_ (.A(_01127_),
    .B(_01131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_2 _19967_ (.A(_01143_),
    .B(_01145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01191_));
 sky130_fd_sc_hd__o211ai_2 _19968_ (.A1(_01127_),
    .A2(_01131_),
    .B1(_01142_),
    .C1(_01191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01193_));
 sky130_fd_sc_hd__and3_2 _19969_ (.A(_01143_),
    .B(_01149_),
    .C(_01190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01194_));
 sky130_fd_sc_hd__nand3_2 _19970_ (.A(_01143_),
    .B(_01149_),
    .C(_01190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01195_));
 sky130_fd_sc_hd__o21ai_2 _19971_ (.A1(_09253_),
    .A2(_09384_),
    .B1(_01193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01196_));
 sky130_fd_sc_hd__o2bb2ai_2 _19972_ (.A1_N(_01193_),
    .A2_N(_01195_),
    .B1(_09253_),
    .B2(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01197_));
 sky130_fd_sc_hd__nand3_2 _19973_ (.A(_01193_),
    .B(\b_l[15] ),
    .C(\a_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01198_));
 sky130_fd_sc_hd__nand4_2 _19974_ (.A(_01195_),
    .B(\a_l[8] ),
    .C(_01193_),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01199_));
 sky130_fd_sc_hd__o21ai_2 _19975_ (.A1(_01194_),
    .A2(_01198_),
    .B1(_01197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01200_));
 sky130_fd_sc_hd__and3_2 _19976_ (.A(_00872_),
    .B(\a_l[15] ),
    .C(\b_l[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01201_));
 sky130_fd_sc_hd__a211o_2 _19977_ (.A1(\b_l[7] ),
    .A2(\a_l[14] ),
    .B1(_09373_),
    .C1(_09264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01202_));
 sky130_fd_sc_hd__nand2_2 _19978_ (.A(\a_l[9] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_2 _19979_ (.A(\a_l[11] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_2 _19980_ (.A(\a_l[10] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01206_));
 sky130_fd_sc_hd__o22a_2 _19981_ (.A1(_09297_),
    .A2(_09329_),
    .B1(_09351_),
    .B2(_09286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01207_));
 sky130_fd_sc_hd__nand2_2 _19982_ (.A(_01205_),
    .B(_01206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01208_));
 sky130_fd_sc_hd__and4_2 _19983_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01209_));
 sky130_fd_sc_hd__nand4_2 _19984_ (.A(\a_l[10] ),
    .B(\a_l[11] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01210_));
 sky130_fd_sc_hd__and3_2 _19985_ (.A(_01210_),
    .B(\b_l[14] ),
    .C(\a_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01211_));
 sky130_fd_sc_hd__and4_2 _19986_ (.A(_01208_),
    .B(_01210_),
    .C(\a_l[9] ),
    .D(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01212_));
 sky130_fd_sc_hd__a22oi_2 _19987_ (.A1(\a_l[9] ),
    .A2(\b_l[14] ),
    .B1(_01208_),
    .B2(_01210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01213_));
 sky130_fd_sc_hd__a21oi_2 _19988_ (.A1(_01211_),
    .A2(_01208_),
    .B1(_01213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01215_));
 sky130_fd_sc_hd__and2_2 _19989_ (.A(\b_l[11] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01216_));
 sky130_fd_sc_hd__nand2_2 _19990_ (.A(\b_l[11] ),
    .B(\a_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_2 _19991_ (.A(\b_l[10] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01218_));
 sky130_fd_sc_hd__nand4_2 _19992_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_l[13] ),
    .D(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_2 _19993_ (.A(\b_l[10] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_2 _19994_ (.A(\b_l[9] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01221_));
 sky130_fd_sc_hd__a22oi_2 _19995_ (.A1(\b_l[10] ),
    .A2(\a_l[13] ),
    .B1(\a_l[14] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_2 _19996_ (.A(_01220_),
    .B(_01221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01223_));
 sky130_fd_sc_hd__o2bb2ai_2 _19997_ (.A1_N(_01220_),
    .A2_N(_01221_),
    .B1(_01110_),
    .B2(_01218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01224_));
 sky130_fd_sc_hd__o221ai_2 _19998_ (.A1(_09308_),
    .A2(_09319_),
    .B1(_01110_),
    .B2(_01218_),
    .C1(_01223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01226_));
 sky130_fd_sc_hd__nand2_2 _19999_ (.A(_01224_),
    .B(_01216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01227_));
 sky130_fd_sc_hd__o2bb2ai_2 _20000_ (.A1_N(_01219_),
    .A2_N(_01223_),
    .B1(_09308_),
    .B2(_09319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01228_));
 sky130_fd_sc_hd__o211ai_2 _20001_ (.A1(_01110_),
    .A2(_01218_),
    .B1(_01216_),
    .C1(_01223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01229_));
 sky130_fd_sc_hd__o22ai_2 _20002_ (.A1(_09340_),
    .A2(_01111_),
    .B1(_01109_),
    .B2(_01113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_2 _20003_ (.A(_01114_),
    .B(_01122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01231_));
 sky130_fd_sc_hd__nand3_2 _20004_ (.A(_01226_),
    .B(_01227_),
    .C(_01231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01232_));
 sky130_fd_sc_hd__nand3_2 _20005_ (.A(_01228_),
    .B(_01229_),
    .C(_01230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01233_));
 sky130_fd_sc_hd__inv_2 _20006_ (.A(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01234_));
 sky130_fd_sc_hd__and3_2 _20007_ (.A(_01215_),
    .B(_01232_),
    .C(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01235_));
 sky130_fd_sc_hd__nand3_2 _20008_ (.A(_01215_),
    .B(_01232_),
    .C(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01237_));
 sky130_fd_sc_hd__a21oi_2 _20009_ (.A1(_01232_),
    .A2(_01233_),
    .B1(_01215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01238_));
 sky130_fd_sc_hd__a21o_2 _20010_ (.A1(_01232_),
    .A2(_01233_),
    .B1(_01215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01239_));
 sky130_fd_sc_hd__nand2_2 _20011_ (.A(_01237_),
    .B(_01239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01240_));
 sky130_fd_sc_hd__a22oi_2 _20012_ (.A1(_01103_),
    .A2(_01099_),
    .B1(_01239_),
    .B2(_01237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01241_));
 sky130_fd_sc_hd__o22ai_2 _20013_ (.A1(_01104_),
    .A2(_01098_),
    .B1(_01238_),
    .B2(_01235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01242_));
 sky130_fd_sc_hd__nor3_2 _20014_ (.A(_01238_),
    .B(_01105_),
    .C(_01235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01243_));
 sky130_fd_sc_hd__nand4_2 _20015_ (.A(_01099_),
    .B(_01239_),
    .C(_01103_),
    .D(_01237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01244_));
 sky130_fd_sc_hd__a21o_2 _20016_ (.A1(_01124_),
    .A2(_01134_),
    .B1(_01121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01245_));
 sky130_fd_sc_hd__o21bai_2 _20017_ (.A1(_01241_),
    .A2(_01243_),
    .B1_N(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01246_));
 sky130_fd_sc_hd__a22oi_2 _20018_ (.A1(_01120_),
    .A2(_01136_),
    .B1(_01240_),
    .B2(_01105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01247_));
 sky130_fd_sc_hd__nand3_2 _20019_ (.A(_01242_),
    .B(_01244_),
    .C(_01245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01248_));
 sky130_fd_sc_hd__nand4_2 _20020_ (.A(_01120_),
    .B(_01136_),
    .C(_01242_),
    .D(_01244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01249_));
 sky130_fd_sc_hd__o22ai_2 _20021_ (.A1(_01121_),
    .A2(_01137_),
    .B1(_01241_),
    .B2(_01243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01250_));
 sky130_fd_sc_hd__nand3_2 _20022_ (.A(_01202_),
    .B(_01249_),
    .C(_01250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01251_));
 sky130_fd_sc_hd__nand3_2 _20023_ (.A(_01246_),
    .B(_01248_),
    .C(_01201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01252_));
 sky130_fd_sc_hd__nand2_2 _20024_ (.A(_01251_),
    .B(_01252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01253_));
 sky130_fd_sc_hd__nand3_2 _20025_ (.A(_01152_),
    .B(_01251_),
    .C(_01252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01254_));
 sky130_fd_sc_hd__a21oi_2 _20026_ (.A1(_01251_),
    .A2(_01252_),
    .B1(_01152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_2 _20027_ (.A(_01153_),
    .B(_01253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01256_));
 sky130_fd_sc_hd__nand3_2 _20028_ (.A(_01256_),
    .B(_01200_),
    .C(_01254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01258_));
 sky130_fd_sc_hd__a21o_2 _20029_ (.A1(_01254_),
    .A2(_01256_),
    .B1(_01200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01259_));
 sky130_fd_sc_hd__a22o_2 _20030_ (.A1(_01197_),
    .A2(_01199_),
    .B1(_01254_),
    .B2(_01256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01260_));
 sky130_fd_sc_hd__o2111ai_2 _20031_ (.A1(_01198_),
    .A2(_01194_),
    .B1(_01197_),
    .C1(_01254_),
    .D1(_01256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01261_));
 sky130_fd_sc_hd__o211ai_2 _20032_ (.A1(_01159_),
    .A2(_01188_),
    .B1(_01258_),
    .C1(_01259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01262_));
 sky130_fd_sc_hd__nand3_2 _20033_ (.A(_01189_),
    .B(_01260_),
    .C(_01261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01263_));
 sky130_fd_sc_hd__nand2_2 _20034_ (.A(_01262_),
    .B(_01263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01264_));
 sky130_fd_sc_hd__o31ai_2 _20035_ (.A1(_09242_),
    .A2(_09384_),
    .A3(_01092_),
    .B1(_01090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01265_));
 sky130_fd_sc_hd__nand3_2 _20036_ (.A(_01262_),
    .B(_01263_),
    .C(_01265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01266_));
 sky130_fd_sc_hd__a21o_2 _20037_ (.A1(_01262_),
    .A2(_01263_),
    .B1(_01265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01267_));
 sky130_fd_sc_hd__o2111ai_2 _20038_ (.A1(_01086_),
    .A2(_01165_),
    .B1(_01175_),
    .C1(_01266_),
    .D1(_01267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_2 _20039_ (.A(_01265_),
    .B(_01264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01270_));
 sky130_fd_sc_hd__o2bb2ai_2 _20040_ (.A1_N(_01265_),
    .A2_N(_01264_),
    .B1(_01174_),
    .B2(_01167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_2 _20041_ (.A(_01270_),
    .B(_01271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01272_));
 sky130_fd_sc_hd__o21a_2 _20042_ (.A1(_01270_),
    .A2(_01271_),
    .B1(_01269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01273_));
 sky130_fd_sc_hd__o21ai_2 _20043_ (.A1(_01270_),
    .A2(_01271_),
    .B1(_01269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01274_));
 sky130_fd_sc_hd__a21oi_2 _20044_ (.A1(_01179_),
    .A2(_01187_),
    .B1(_01274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01275_));
 sky130_fd_sc_hd__a31o_2 _20045_ (.A1(_01179_),
    .A2(_01187_),
    .A3(_01274_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01276_));
 sky130_fd_sc_hd__nor2_2 _20046_ (.A(_01275_),
    .B(_01276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00393_));
 sky130_fd_sc_hd__a31o_2 _20047_ (.A1(_01189_),
    .A2(_01260_),
    .A3(_01261_),
    .B1(_01265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01277_));
 sky130_fd_sc_hd__o21ai_2 _20048_ (.A1(_01200_),
    .A2(_01255_),
    .B1(_01254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01279_));
 sky130_fd_sc_hd__o21a_2 _20049_ (.A1(_01200_),
    .A2(_01255_),
    .B1(_01254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_2 _20050_ (.A(\a_l[11] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_2 _20051_ (.A(\a_l[12] ),
    .B(\b_l[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_2 _20052_ (.A(\a_l[12] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01283_));
 sky130_fd_sc_hd__and4_2 _20053_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01284_));
 sky130_fd_sc_hd__nand4_2 _20054_ (.A(\a_l[11] ),
    .B(\a_l[12] ),
    .C(\b_l[12] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_2 _20055_ (.A(_01281_),
    .B(_01282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01286_));
 sky130_fd_sc_hd__and4_2 _20056_ (.A(_01286_),
    .B(\b_l[14] ),
    .C(\a_l[10] ),
    .D(_01285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01287_));
 sky130_fd_sc_hd__o2111ai_2 _20057_ (.A1(_01205_),
    .A2(_01283_),
    .B1(\a_l[10] ),
    .C1(\b_l[14] ),
    .D1(_01286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01288_));
 sky130_fd_sc_hd__o2bb2a_2 _20058_ (.A1_N(_01285_),
    .A2_N(_01286_),
    .B1(_09286_),
    .B2(_09362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01290_));
 sky130_fd_sc_hd__a22o_2 _20059_ (.A1(\a_l[10] ),
    .A2(\b_l[14] ),
    .B1(_01285_),
    .B2(_01286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01291_));
 sky130_fd_sc_hd__nand2_2 _20060_ (.A(_01288_),
    .B(_01291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_2 _20061_ (.A(\b_l[11] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_2 _20062_ (.A(\b_l[10] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01294_));
 sky130_fd_sc_hd__nand4_2 _20063_ (.A(\b_l[9] ),
    .B(\b_l[10] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_2 _20064_ (.A(\b_l[9] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01296_));
 sky130_fd_sc_hd__a22oi_2 _20065_ (.A1(\b_l[10] ),
    .A2(\a_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_2 _20066_ (.A(_01218_),
    .B(_01296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01298_));
 sky130_fd_sc_hd__o2bb2ai_2 _20067_ (.A1_N(_01295_),
    .A2_N(_01298_),
    .B1(_09308_),
    .B2(_09340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01299_));
 sky130_fd_sc_hd__a41o_2 _20068_ (.A1(\b_l[9] ),
    .A2(\b_l[10] ),
    .A3(\a_l[14] ),
    .A4(\a_l[15] ),
    .B1(_01293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01301_));
 sky130_fd_sc_hd__o2111ai_2 _20069_ (.A1(_01221_),
    .A2(_01294_),
    .B1(\b_l[11] ),
    .C1(\a_l[13] ),
    .D1(_01298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01302_));
 sky130_fd_sc_hd__o22a_2 _20070_ (.A1(_09308_),
    .A2(_09319_),
    .B1(_01110_),
    .B2(_01218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01303_));
 sky130_fd_sc_hd__o21ai_2 _20071_ (.A1(_01217_),
    .A2(_01222_),
    .B1(_01219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01304_));
 sky130_fd_sc_hd__o211a_2 _20072_ (.A1(_01297_),
    .A2(_01301_),
    .B1(_01304_),
    .C1(_01299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01305_));
 sky130_fd_sc_hd__o211ai_2 _20073_ (.A1(_01297_),
    .A2(_01301_),
    .B1(_01304_),
    .C1(_01299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01306_));
 sky130_fd_sc_hd__a21oi_2 _20074_ (.A1(_01299_),
    .A2(_01302_),
    .B1(_01304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01307_));
 sky130_fd_sc_hd__o2bb2ai_2 _20075_ (.A1_N(_01299_),
    .A2_N(_01302_),
    .B1(_01303_),
    .B2(_01222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01308_));
 sky130_fd_sc_hd__a21oi_2 _20076_ (.A1(_01306_),
    .A2(_01308_),
    .B1(_01292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01309_));
 sky130_fd_sc_hd__o211ai_2 _20077_ (.A1(_01287_),
    .A2(_01290_),
    .B1(_01306_),
    .C1(_01308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01310_));
 sky130_fd_sc_hd__o22ai_2 _20078_ (.A1(_01287_),
    .A2(_01290_),
    .B1(_01305_),
    .B2(_01307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01312_));
 sky130_fd_sc_hd__nand3b_2 _20079_ (.A_N(_01292_),
    .B(_01306_),
    .C(_01308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01313_));
 sky130_fd_sc_hd__o21ai_2 _20080_ (.A1(_00872_),
    .A2(_01100_),
    .B1(_01310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01314_));
 sky130_fd_sc_hd__a21o_2 _20081_ (.A1(_01312_),
    .A2(_01313_),
    .B1(_01101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01315_));
 sky130_fd_sc_hd__nand3_2 _20082_ (.A(_01312_),
    .B(_01313_),
    .C(_01101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01316_));
 sky130_fd_sc_hd__a311oi_2 _20083_ (.A1(_01226_),
    .A2(_01227_),
    .A3(_01231_),
    .B1(_01213_),
    .C1(_01212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01317_));
 sky130_fd_sc_hd__a21bo_2 _20084_ (.A1(_01215_),
    .A2(_01232_),
    .B1_N(_01233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01318_));
 sky130_fd_sc_hd__a21o_2 _20085_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01319_));
 sky130_fd_sc_hd__o221ai_2 _20086_ (.A1(_01234_),
    .A2(_01317_),
    .B1(_01309_),
    .B2(_01314_),
    .C1(_01316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01320_));
 sky130_fd_sc_hd__a32o_2 _20087_ (.A1(_01201_),
    .A2(_01246_),
    .A3(_01248_),
    .B1(_01319_),
    .B2(_01320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01321_));
 sky130_fd_sc_hd__nand3b_2 _20088_ (.A_N(_01252_),
    .B(_01319_),
    .C(_01320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01323_));
 sky130_fd_sc_hd__nand2_2 _20089_ (.A(_01321_),
    .B(_01323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_2 _20090_ (.A(\a_l[9] ),
    .B(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01325_));
 sky130_fd_sc_hd__o22ai_2 _20091_ (.A1(_01209_),
    .A2(_01212_),
    .B1(_01243_),
    .B2(_01247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01326_));
 sky130_fd_sc_hd__o2111ai_2 _20092_ (.A1(_01204_),
    .A2(_01207_),
    .B1(_01210_),
    .C1(_01244_),
    .D1(_01248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_2 _20093_ (.A(_01326_),
    .B(_01327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01328_));
 sky130_fd_sc_hd__a21o_2 _20094_ (.A1(_01326_),
    .A2(_01327_),
    .B1(_01325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01329_));
 sky130_fd_sc_hd__o211ai_2 _20095_ (.A1(_09275_),
    .A2(_09384_),
    .B1(_01326_),
    .C1(_01327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_2 _20096_ (.A(_01329_),
    .B(_01330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01331_));
 sky130_fd_sc_hd__nand3_2 _20097_ (.A(_01323_),
    .B(_01329_),
    .C(_01330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01332_));
 sky130_fd_sc_hd__nand4_2 _20098_ (.A(_01321_),
    .B(_01323_),
    .C(_01329_),
    .D(_01330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_2 _20099_ (.A(_01324_),
    .B(_01331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01335_));
 sky130_fd_sc_hd__nand3_2 _20100_ (.A(_01331_),
    .B(_01323_),
    .C(_01321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01336_));
 sky130_fd_sc_hd__nand3_2 _20101_ (.A(_01324_),
    .B(_01329_),
    .C(_01330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01337_));
 sky130_fd_sc_hd__nand3_2 _20102_ (.A(_01280_),
    .B(_01334_),
    .C(_01335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01338_));
 sky130_fd_sc_hd__nand3_2 _20103_ (.A(_01337_),
    .B(_01279_),
    .C(_01336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01339_));
 sky130_fd_sc_hd__a22o_2 _20104_ (.A1(_01195_),
    .A2(_01196_),
    .B1(_01338_),
    .B2(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01340_));
 sky130_fd_sc_hd__nand4_2 _20105_ (.A(_01195_),
    .B(_01196_),
    .C(_01338_),
    .D(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01341_));
 sky130_fd_sc_hd__o311ai_2 _20106_ (.A1(_09253_),
    .A2(_01194_),
    .A3(_09384_),
    .B1(_01193_),
    .C1(_01339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01342_));
 sky130_fd_sc_hd__a22oi_2 _20107_ (.A1(_01262_),
    .A2(_01277_),
    .B1(_01340_),
    .B2(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01343_));
 sky130_fd_sc_hd__nand4_2 _20108_ (.A(_01262_),
    .B(_01277_),
    .C(_01340_),
    .D(_01341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2b_2 _20109_ (.A_N(_01343_),
    .B(_01344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01345_));
 sky130_fd_sc_hd__o2111ai_2 _20110_ (.A1(_01270_),
    .A2(_01271_),
    .B1(_01179_),
    .C1(_01181_),
    .D1(_01269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01346_));
 sky130_fd_sc_hd__nand3_2 _20111_ (.A(_01182_),
    .B(_01183_),
    .C(_01273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01347_));
 sky130_fd_sc_hd__o21a_2 _20112_ (.A1(_01179_),
    .A2(_01272_),
    .B1(_01269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01348_));
 sky130_fd_sc_hd__o211a_2 _20113_ (.A1(_01272_),
    .A2(_01179_),
    .B1(_01269_),
    .C1(_01347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01349_));
 sky130_fd_sc_hd__nand3_2 _20114_ (.A(_00975_),
    .B(_00976_),
    .C(_01349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01350_));
 sky130_fd_sc_hd__o211ai_2 _20115_ (.A1(_01184_),
    .A2(_01346_),
    .B1(_01348_),
    .C1(_01347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_2 _20116_ (.A(_01350_),
    .B(_01351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_2 _20117_ (.A(_01352_),
    .B(_01345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01353_));
 sky130_fd_sc_hd__nand3b_2 _20118_ (.A_N(_01345_),
    .B(_01350_),
    .C(_01351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01355_));
 sky130_fd_sc_hd__and3_2 _20119_ (.A(_09690_),
    .B(_01353_),
    .C(_01355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00394_));
 sky130_fd_sc_hd__o31a_2 _20120_ (.A1(_09275_),
    .A2(_09384_),
    .A3(_01328_),
    .B1(_01326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01356_));
 sky130_fd_sc_hd__inv_2 _20121_ (.A(_01356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01357_));
 sky130_fd_sc_hd__o21ai_2 _20122_ (.A1(_01292_),
    .A2(_01307_),
    .B1(_01306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01358_));
 sky130_fd_sc_hd__o21ai_2 _20123_ (.A1(_01293_),
    .A2(_01297_),
    .B1(_01295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_2 _20124_ (.A(\b_l[11] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_2 _20125_ (.A(\b_l[11] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01361_));
 sky130_fd_sc_hd__nand2_2 _20126_ (.A(_01294_),
    .B(_01360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01362_));
 sky130_fd_sc_hd__o21a_2 _20127_ (.A1(_01218_),
    .A2(_01361_),
    .B1(_01362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01363_));
 sky130_fd_sc_hd__o21ai_2 _20128_ (.A1(_01218_),
    .A2(_01361_),
    .B1(_01362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_2 _20129_ (.A(_01359_),
    .B(_01363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01366_));
 sky130_fd_sc_hd__o211ai_2 _20130_ (.A1(_01297_),
    .A2(_01293_),
    .B1(_01295_),
    .C1(_01365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01367_));
 sky130_fd_sc_hd__and2_2 _20131_ (.A(\a_l[11] ),
    .B(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_2 _20132_ (.A(\b_l[12] ),
    .B(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01369_));
 sky130_fd_sc_hd__nand3_2 _20133_ (.A(\a_l[12] ),
    .B(\b_l[12] ),
    .C(\a_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01370_));
 sky130_fd_sc_hd__nand4_2 _20134_ (.A(\a_l[12] ),
    .B(\b_l[12] ),
    .C(\a_l[13] ),
    .D(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2_2 _20135_ (.A(_01283_),
    .B(_01369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01372_));
 sky130_fd_sc_hd__a2bb2oi_2 _20136_ (.A1_N(_09297_),
    .A2_N(_09362_),
    .B1(_01371_),
    .B2(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01373_));
 sky130_fd_sc_hd__a22o_2 _20137_ (.A1(\a_l[11] ),
    .A2(\b_l[14] ),
    .B1(_01371_),
    .B2(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01374_));
 sky130_fd_sc_hd__o211a_2 _20138_ (.A1(_09351_),
    .A2(_01370_),
    .B1(_01368_),
    .C1(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01376_));
 sky130_fd_sc_hd__o2111ai_2 _20139_ (.A1(_09351_),
    .A2(_01370_),
    .B1(\b_l[14] ),
    .C1(\a_l[11] ),
    .D1(_01372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01377_));
 sky130_fd_sc_hd__a22o_2 _20140_ (.A1(_01366_),
    .A2(_01367_),
    .B1(_01374_),
    .B2(_01377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01378_));
 sky130_fd_sc_hd__nand4_2 _20141_ (.A(_01366_),
    .B(_01367_),
    .C(_01374_),
    .D(_01377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_2 _20142_ (.A(_01378_),
    .B(_01379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01380_));
 sky130_fd_sc_hd__xnor2_2 _20143_ (.A(_01358_),
    .B(_01380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01381_));
 sky130_fd_sc_hd__o31a_2 _20144_ (.A1(_09319_),
    .A2(_09351_),
    .A3(_01205_),
    .B1(_01288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01382_));
 sky130_fd_sc_hd__a31o_2 _20145_ (.A1(_01312_),
    .A2(_01313_),
    .A3(_01101_),
    .B1(_01318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01383_));
 sky130_fd_sc_hd__o22ai_2 _20146_ (.A1(_01234_),
    .A2(_01317_),
    .B1(_01309_),
    .B2(_01314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01384_));
 sky130_fd_sc_hd__and3_2 _20147_ (.A(_01316_),
    .B(_01384_),
    .C(_01382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01385_));
 sky130_fd_sc_hd__nand3_2 _20148_ (.A(_01316_),
    .B(_01384_),
    .C(_01382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01387_));
 sky130_fd_sc_hd__o211ai_2 _20149_ (.A1(_01284_),
    .A2(_01287_),
    .B1(_01315_),
    .C1(_01383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01388_));
 sky130_fd_sc_hd__nand4_2 _20150_ (.A(_01388_),
    .B(\a_l[10] ),
    .C(_01387_),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01389_));
 sky130_fd_sc_hd__o2bb2ai_2 _20151_ (.A1_N(_01387_),
    .A2_N(_01388_),
    .B1(_09286_),
    .B2(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01390_));
 sky130_fd_sc_hd__a21oi_2 _20152_ (.A1(_01389_),
    .A2(_01390_),
    .B1(_01381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01391_));
 sky130_fd_sc_hd__a21o_2 _20153_ (.A1(_01389_),
    .A2(_01390_),
    .B1(_01381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01392_));
 sky130_fd_sc_hd__nand3_2 _20154_ (.A(_01390_),
    .B(_01381_),
    .C(_01389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01393_));
 sky130_fd_sc_hd__inv_2 _20155_ (.A(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01394_));
 sky130_fd_sc_hd__o2bb2ai_2 _20156_ (.A1_N(_01321_),
    .A2_N(_01332_),
    .B1(_01391_),
    .B2(_01394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01395_));
 sky130_fd_sc_hd__nand4_2 _20157_ (.A(_01321_),
    .B(_01332_),
    .C(_01392_),
    .D(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_2 _20158_ (.A(_01357_),
    .B(_01395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01398_));
 sky130_fd_sc_hd__a41o_2 _20159_ (.A1(_01321_),
    .A2(_01332_),
    .A3(_01392_),
    .A4(_01393_),
    .B1(_01398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01399_));
 sky130_fd_sc_hd__a21o_2 _20160_ (.A1(_01395_),
    .A2(_01396_),
    .B1(_01357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01400_));
 sky130_fd_sc_hd__a22oi_2 _20161_ (.A1(_01338_),
    .A2(_01342_),
    .B1(_01399_),
    .B2(_01400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01401_));
 sky130_fd_sc_hd__a22o_2 _20162_ (.A1(_01338_),
    .A2(_01342_),
    .B1(_01399_),
    .B2(_01400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01402_));
 sky130_fd_sc_hd__nand4_2 _20163_ (.A(_01338_),
    .B(_01342_),
    .C(_01399_),
    .D(_01400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01403_));
 sky130_fd_sc_hd__nand2_2 _20164_ (.A(_01402_),
    .B(_01403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01404_));
 sky130_fd_sc_hd__a21o_2 _20165_ (.A1(_01344_),
    .A2(_01355_),
    .B1(_01404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01405_));
 sky130_fd_sc_hd__o211ai_2 _20166_ (.A1(_01345_),
    .A2(_01352_),
    .B1(_01404_),
    .C1(_01344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01406_));
 sky130_fd_sc_hd__and3_2 _20167_ (.A(_09690_),
    .B(_01405_),
    .C(_01406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00395_));
 sky130_fd_sc_hd__o31ai_2 _20168_ (.A1(_09286_),
    .A2(_09384_),
    .A3(_01385_),
    .B1(_01388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01407_));
 sky130_fd_sc_hd__a21o_2 _20169_ (.A1(\b_l[10] ),
    .A2(\a_l[14] ),
    .B1(_09308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01408_));
 sky130_fd_sc_hd__and3_2 _20170_ (.A(_01218_),
    .B(\a_l[15] ),
    .C(\b_l[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01409_));
 sky130_fd_sc_hd__nand2_2 _20171_ (.A(\b_l[13] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_2 _20172_ (.A(\a_l[13] ),
    .B(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_2 _20173_ (.A(\b_l[12] ),
    .B(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01412_));
 sky130_fd_sc_hd__nand4_2 _20174_ (.A(\b_l[12] ),
    .B(\a_l[13] ),
    .C(\b_l[13] ),
    .D(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01413_));
 sky130_fd_sc_hd__nand2_2 _20175_ (.A(_01411_),
    .B(_01412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01414_));
 sky130_fd_sc_hd__o2bb2ai_2 _20176_ (.A1_N(_01413_),
    .A2_N(_01414_),
    .B1(_09319_),
    .B2(_09362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01415_));
 sky130_fd_sc_hd__o2111ai_2 _20177_ (.A1(_01369_),
    .A2(_01410_),
    .B1(\a_l[12] ),
    .C1(\b_l[14] ),
    .D1(_01414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01416_));
 sky130_fd_sc_hd__o2bb2ai_2 _20178_ (.A1_N(_01415_),
    .A2_N(_01416_),
    .B1(_09373_),
    .B2(_01408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01418_));
 sky130_fd_sc_hd__nand3_2 _20179_ (.A(_01415_),
    .B(_01416_),
    .C(_01409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01419_));
 sky130_fd_sc_hd__o2bb2ai_2 _20180_ (.A1_N(_01359_),
    .A2_N(_01363_),
    .B1(_01373_),
    .B2(_01376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01420_));
 sky130_fd_sc_hd__nand3_2 _20181_ (.A(_01367_),
    .B(_01374_),
    .C(_01377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01421_));
 sky130_fd_sc_hd__nand2_2 _20182_ (.A(_01366_),
    .B(_01421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01422_));
 sky130_fd_sc_hd__a21oi_2 _20183_ (.A1(_01418_),
    .A2(_01419_),
    .B1(_01422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01423_));
 sky130_fd_sc_hd__nand4_2 _20184_ (.A(_01367_),
    .B(_01418_),
    .C(_01419_),
    .D(_01420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01424_));
 sky130_fd_sc_hd__and2b_2 _20185_ (.A_N(_01423_),
    .B(_01424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01425_));
 sky130_fd_sc_hd__nor2_2 _20186_ (.A(_09297_),
    .B(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01426_));
 sky130_fd_sc_hd__a41o_2 _20187_ (.A1(\a_l[12] ),
    .A2(\b_l[12] ),
    .A3(\a_l[13] ),
    .A4(\b_l[13] ),
    .B1(_01376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01427_));
 sky130_fd_sc_hd__a31oi_2 _20188_ (.A1(_01358_),
    .A2(_01378_),
    .A3(_01379_),
    .B1(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01429_));
 sky130_fd_sc_hd__a31o_2 _20189_ (.A1(_01358_),
    .A2(_01378_),
    .A3(_01379_),
    .B1(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01430_));
 sky130_fd_sc_hd__nand4_2 _20190_ (.A(_01358_),
    .B(_01378_),
    .C(_01379_),
    .D(_01427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_2 _20191_ (.A(_01431_),
    .B(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01432_));
 sky130_fd_sc_hd__and3_2 _20192_ (.A(_01430_),
    .B(_01431_),
    .C(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01433_));
 sky130_fd_sc_hd__a21oi_2 _20193_ (.A1(_01430_),
    .A2(_01431_),
    .B1(_01426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01434_));
 sky130_fd_sc_hd__o21ba_2 _20194_ (.A1(_01433_),
    .A2(_01434_),
    .B1_N(_01425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01435_));
 sky130_fd_sc_hd__o21ai_2 _20195_ (.A1(_01429_),
    .A2(_01432_),
    .B1(_01425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_2 _20196_ (.A(_01434_),
    .B(_01436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01437_));
 sky130_fd_sc_hd__o21a_2 _20197_ (.A1(_01435_),
    .A2(_01437_),
    .B1(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01438_));
 sky130_fd_sc_hd__o21ai_2 _20198_ (.A1(_01435_),
    .A2(_01437_),
    .B1(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01440_));
 sky130_fd_sc_hd__nor3_2 _20199_ (.A(_01435_),
    .B(_01437_),
    .C(_01393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_2 _20200_ (.A(_01440_),
    .B(_01407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_2 _20201_ (.A(_01441_),
    .B(_01442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01443_));
 sky130_fd_sc_hd__o21bai_2 _20202_ (.A1(_01438_),
    .A2(_01441_),
    .B1_N(_01407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01444_));
 sky130_fd_sc_hd__o21ai_2 _20203_ (.A1(_01441_),
    .A2(_01442_),
    .B1(_01444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01445_));
 sky130_fd_sc_hd__a21bo_2 _20204_ (.A1(_01396_),
    .A2(_01398_),
    .B1_N(_01444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01446_));
 sky130_fd_sc_hd__a21oi_2 _20205_ (.A1(_01396_),
    .A2(_01398_),
    .B1(_01445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01447_));
 sky130_fd_sc_hd__a21o_2 _20206_ (.A1(_01396_),
    .A2(_01398_),
    .B1(_01445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01448_));
 sky130_fd_sc_hd__nand3_2 _20207_ (.A(_01396_),
    .B(_01398_),
    .C(_01445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01449_));
 sky130_fd_sc_hd__o21ai_2 _20208_ (.A1(_01443_),
    .A2(_01446_),
    .B1(_01449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01451_));
 sky130_fd_sc_hd__and4b_2 _20209_ (.A_N(_01343_),
    .B(_01344_),
    .C(_01402_),
    .D(_01403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01452_));
 sky130_fd_sc_hd__and2_2 _20210_ (.A(_01351_),
    .B(_01452_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01453_));
 sky130_fd_sc_hd__o21ai_2 _20211_ (.A1(_01344_),
    .A2(_01401_),
    .B1(_01403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01454_));
 sky130_fd_sc_hd__a21oi_2 _20212_ (.A1(_01350_),
    .A2(_01453_),
    .B1(_01454_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01455_));
 sky130_fd_sc_hd__o21ai_2 _20213_ (.A1(_01451_),
    .A2(_01455_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01456_));
 sky130_fd_sc_hd__a21oi_2 _20214_ (.A1(_01451_),
    .A2(_01455_),
    .B1(_01456_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00396_));
 sky130_fd_sc_hd__a21o_2 _20215_ (.A1(_01440_),
    .A2(_01407_),
    .B1(_01441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01457_));
 sky130_fd_sc_hd__o21ai_2 _20216_ (.A1(_01218_),
    .A2(_01361_),
    .B1(_01419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_2 _20217_ (.A(\b_l[12] ),
    .B(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_2 _20218_ (.A(_01410_),
    .B(_01459_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01461_));
 sky130_fd_sc_hd__nand4_2 _20219_ (.A(\b_l[12] ),
    .B(\b_l[13] ),
    .C(\a_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01462_));
 sky130_fd_sc_hd__nand4_2 _20220_ (.A(_01461_),
    .B(_01462_),
    .C(\a_l[13] ),
    .D(\b_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01463_));
 sky130_fd_sc_hd__o2bb2ai_2 _20221_ (.A1_N(_01461_),
    .A2_N(_01462_),
    .B1(_09340_),
    .B2(_09362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01464_));
 sky130_fd_sc_hd__and2_2 _20222_ (.A(_01463_),
    .B(_01464_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_2 _20223_ (.A(_01458_),
    .B(_01465_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01466_));
 sky130_fd_sc_hd__or2_2 _20224_ (.A(_01465_),
    .B(_01458_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01467_));
 sky130_fd_sc_hd__nand2_2 _20225_ (.A(_01466_),
    .B(_01467_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_2 _20226_ (.A(_09319_),
    .B(_09384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01469_));
 sky130_fd_sc_hd__o21ai_2 _20227_ (.A1(_01411_),
    .A2(_01412_),
    .B1(_01416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01470_));
 sky130_fd_sc_hd__o211ai_2 _20228_ (.A1(_01369_),
    .A2(_01410_),
    .B1(_01416_),
    .C1(_01424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01472_));
 sky130_fd_sc_hd__nand4_2 _20229_ (.A(_01422_),
    .B(_01470_),
    .C(_01418_),
    .D(_01419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01473_));
 sky130_fd_sc_hd__a21oi_2 _20230_ (.A1(_01472_),
    .A2(_01473_),
    .B1(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01474_));
 sky130_fd_sc_hd__a22o_2 _20231_ (.A1(\a_l[12] ),
    .A2(\b_l[15] ),
    .B1(_01472_),
    .B2(_01473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01475_));
 sky130_fd_sc_hd__and3_2 _20232_ (.A(_01472_),
    .B(_01473_),
    .C(_01469_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01476_));
 sky130_fd_sc_hd__o21ai_2 _20233_ (.A1(_01474_),
    .A2(_01476_),
    .B1(_01468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01477_));
 sky130_fd_sc_hd__a31oi_2 _20234_ (.A1(_01469_),
    .A2(_01472_),
    .A3(_01473_),
    .B1(_01468_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_2 _20235_ (.A(_01478_),
    .B(_01475_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01479_));
 sky130_fd_sc_hd__a2bb2o_2 _20236_ (.A1_N(_01436_),
    .A2_N(_01434_),
    .B1(_01479_),
    .B2(_01477_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01480_));
 sky130_fd_sc_hd__nand3_2 _20237_ (.A(_01437_),
    .B(_01477_),
    .C(_01479_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01481_));
 sky130_fd_sc_hd__o31ai_2 _20238_ (.A1(_09297_),
    .A2(_09384_),
    .A3(_01429_),
    .B1(_01431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01483_));
 sky130_fd_sc_hd__a21oi_2 _20239_ (.A1(_01480_),
    .A2(_01481_),
    .B1(_01483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01484_));
 sky130_fd_sc_hd__nand3_2 _20240_ (.A(_01480_),
    .B(_01481_),
    .C(_01483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01485_));
 sky130_fd_sc_hd__and2b_2 _20241_ (.A_N(_01484_),
    .B(_01485_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01486_));
 sky130_fd_sc_hd__and3b_2 _20242_ (.A_N(_01484_),
    .B(_01485_),
    .C(_01457_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01487_));
 sky130_fd_sc_hd__or2_2 _20243_ (.A(_01457_),
    .B(_01486_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01488_));
 sky130_fd_sc_hd__inv_2 _20244_ (.A(_01488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01489_));
 sky130_fd_sc_hd__and2b_2 _20245_ (.A_N(_01487_),
    .B(_01488_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01490_));
 sky130_fd_sc_hd__o22ai_2 _20246_ (.A1(_01443_),
    .A2(_01446_),
    .B1(_01451_),
    .B2(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01491_));
 sky130_fd_sc_hd__o22ai_2 _20247_ (.A1(_01487_),
    .A2(_01489_),
    .B1(_01451_),
    .B2(_01455_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_2 _20248_ (.A(_01491_),
    .B(_01490_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01494_));
 sky130_fd_sc_hd__o211a_2 _20249_ (.A1(_01492_),
    .A2(_01447_),
    .B1(_09690_),
    .C1(_01494_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00397_));
 sky130_fd_sc_hd__and3_2 _20250_ (.A(_01490_),
    .B(_01449_),
    .C(_01448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01495_));
 sky130_fd_sc_hd__nand3_2 _20251_ (.A(_01490_),
    .B(_01449_),
    .C(_01448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01496_));
 sky130_fd_sc_hd__nor3_2 _20252_ (.A(_01345_),
    .B(_01404_),
    .C(_01496_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01497_));
 sky130_fd_sc_hd__and2_2 _20253_ (.A(_01351_),
    .B(_01497_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01498_));
 sky130_fd_sc_hd__nand2_2 _20254_ (.A(_01350_),
    .B(_01498_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01499_));
 sky130_fd_sc_hd__a221oi_2 _20255_ (.A1(_01447_),
    .A2(_01488_),
    .B1(_01495_),
    .B2(_01454_),
    .C1(_01487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01500_));
 sky130_fd_sc_hd__a221o_2 _20256_ (.A1(_01447_),
    .A2(_01488_),
    .B1(_01495_),
    .B2(_01454_),
    .C1(_01487_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01501_));
 sky130_fd_sc_hd__a21oi_2 _20257_ (.A1(_01350_),
    .A2(_01498_),
    .B1(_01501_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01502_));
 sky130_fd_sc_hd__o311a_2 _20258_ (.A1(_09351_),
    .A2(_09373_),
    .A3(_01412_),
    .B1(_01463_),
    .C1(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01503_));
 sky130_fd_sc_hd__a21o_2 _20259_ (.A1(_01462_),
    .A2(_01463_),
    .B1(_01466_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01504_));
 sky130_fd_sc_hd__inv_2 _20260_ (.A(_01504_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01505_));
 sky130_fd_sc_hd__and4b_2 _20261_ (.A_N(_01503_),
    .B(_01504_),
    .C(\a_l[13] ),
    .D(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01506_));
 sky130_fd_sc_hd__o22a_2 _20262_ (.A1(_09340_),
    .A2(_09384_),
    .B1(_01503_),
    .B2(_01505_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01507_));
 sky130_fd_sc_hd__a22o_2 _20263_ (.A1(\a_l[14] ),
    .A2(\b_l[14] ),
    .B1(\a_l[15] ),
    .B2(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01508_));
 sky130_fd_sc_hd__nand4_2 _20264_ (.A(\b_l[13] ),
    .B(\a_l[14] ),
    .C(\b_l[14] ),
    .D(\a_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01509_));
 sky130_fd_sc_hd__a2bb2oi_2 _20265_ (.A1_N(_01506_),
    .A2_N(_01507_),
    .B1(_01508_),
    .B2(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01510_));
 sky130_fd_sc_hd__and4bb_2 _20266_ (.A_N(_01506_),
    .B_N(_01507_),
    .C(_01508_),
    .D(_01509_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01511_));
 sky130_fd_sc_hd__a2bb2o_2 _20267_ (.A1_N(_01510_),
    .A2_N(_01511_),
    .B1(_01475_),
    .B2(_01478_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01512_));
 sky130_fd_sc_hd__or3_2 _20268_ (.A(_01479_),
    .B(_01510_),
    .C(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01514_));
 sky130_fd_sc_hd__a21boi_2 _20269_ (.A1(_01472_),
    .A2(_01469_),
    .B1_N(_01473_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01515_));
 sky130_fd_sc_hd__a21oi_2 _20270_ (.A1(_01512_),
    .A2(_01514_),
    .B1(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01516_));
 sky130_fd_sc_hd__o31a_2 _20271_ (.A1(_01479_),
    .A2(_01510_),
    .A3(_01511_),
    .B1(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01517_));
 sky130_fd_sc_hd__nand2_2 _20272_ (.A(_01514_),
    .B(_01515_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01518_));
 sky130_fd_sc_hd__a21o_2 _20273_ (.A1(_01512_),
    .A2(_01517_),
    .B1(_01516_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01519_));
 sky130_fd_sc_hd__a32oi_2 _20274_ (.A1(_01437_),
    .A2(_01477_),
    .A3(_01479_),
    .B1(_01480_),
    .B2(_01483_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01520_));
 sky130_fd_sc_hd__and2b_2 _20275_ (.A_N(_01520_),
    .B(_01519_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01521_));
 sky130_fd_sc_hd__nand2_2 _20276_ (.A(_01519_),
    .B(_01520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01522_));
 sky130_fd_sc_hd__or2_2 _20277_ (.A(_01519_),
    .B(_01520_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01523_));
 sky130_fd_sc_hd__and2_2 _20278_ (.A(_01522_),
    .B(_01523_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01525_));
 sky130_fd_sc_hd__a22oi_2 _20279_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01499_),
    .B2(_01500_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01526_));
 sky130_fd_sc_hd__o21ai_2 _20280_ (.A1(_01525_),
    .A2(_01502_),
    .B1(_09690_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01527_));
 sky130_fd_sc_hd__a21oi_2 _20281_ (.A1(_01502_),
    .A2(_01525_),
    .B1(_01527_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_2 _20282_ (.A(\a_l[14] ),
    .B(\b_l[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01528_));
 sky130_fd_sc_hd__o22a_2 _20283_ (.A1(\b_l[15] ),
    .A2(_01410_),
    .B1(_01528_),
    .B2(\b_l[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01529_));
 sky130_fd_sc_hd__or3_2 _20284_ (.A(_09362_),
    .B(_09373_),
    .C(_01529_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01530_));
 sky130_fd_sc_hd__a22o_2 _20285_ (.A1(\b_l[14] ),
    .A2(\a_l[15] ),
    .B1(\b_l[15] ),
    .B2(\a_l[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01531_));
 sky130_fd_sc_hd__o311a_2 _20286_ (.A1(_09362_),
    .A2(_09373_),
    .A3(_01529_),
    .B1(_01531_),
    .C1(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01532_));
 sky130_fd_sc_hd__a21oi_2 _20287_ (.A1(_01530_),
    .A2(_01531_),
    .B1(_01511_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01533_));
 sky130_fd_sc_hd__nor2_2 _20288_ (.A(_01532_),
    .B(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01535_));
 sky130_fd_sc_hd__o21a_2 _20289_ (.A1(_01505_),
    .A2(_01506_),
    .B1(_01535_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01536_));
 sky130_fd_sc_hd__o22a_2 _20290_ (.A1(_01505_),
    .A2(_01506_),
    .B1(_01532_),
    .B2(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01537_));
 sky130_fd_sc_hd__nor4_2 _20291_ (.A(_01505_),
    .B(_01506_),
    .C(_01532_),
    .D(_01533_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01538_));
 sky130_fd_sc_hd__o211a_2 _20292_ (.A1(_01537_),
    .A2(_01538_),
    .B1(_01512_),
    .C1(_01518_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01539_));
 sky130_fd_sc_hd__a211oi_2 _20293_ (.A1(_01512_),
    .A2(_01518_),
    .B1(_01537_),
    .C1(_01538_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01540_));
 sky130_fd_sc_hd__or2_2 _20294_ (.A(_01539_),
    .B(_01540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01541_));
 sky130_fd_sc_hd__o22ai_2 _20295_ (.A1(_01539_),
    .A2(_01540_),
    .B1(_01525_),
    .B2(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01542_));
 sky130_fd_sc_hd__o21bai_2 _20296_ (.A1(_01521_),
    .A2(_01526_),
    .B1_N(_01541_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01543_));
 sky130_fd_sc_hd__o211a_2 _20297_ (.A1(_01542_),
    .A2(_01521_),
    .B1(_09690_),
    .C1(_01543_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00399_));
 sky130_fd_sc_hd__o21a_2 _20298_ (.A1(_09373_),
    .A2(_09384_),
    .B1(_01530_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01544_));
 sky130_fd_sc_hd__a41o_2 _20299_ (.A1(\a_l[14] ),
    .A2(\b_l[14] ),
    .A3(\a_l[15] ),
    .A4(\b_l[15] ),
    .B1(_01544_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01545_));
 sky130_fd_sc_hd__o21ba_2 _20300_ (.A1(_01532_),
    .A2(_01536_),
    .B1_N(_01545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01546_));
 sky130_fd_sc_hd__nor3b_2 _20301_ (.A(_01532_),
    .B(_01536_),
    .C_N(_01545_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_2 _20302_ (.A(_01546_),
    .B(_01547_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_2 _20303_ (.A(_01521_),
    .B(_01539_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_2 _20304_ (.A(_01540_),
    .B(_01549_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01550_));
 sky130_fd_sc_hd__a211o_2 _20305_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01539_),
    .C1(_01540_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_01551_));
 sky130_fd_sc_hd__o22ai_2 _20306_ (.A1(_01540_),
    .A2(_01549_),
    .B1(_01551_),
    .B2(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01552_));
 sky130_fd_sc_hd__o22ai_2 _20307_ (.A1(_01546_),
    .A2(_01547_),
    .B1(_01551_),
    .B2(_01502_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_2 _20308_ (.A(_01552_),
    .B(_01548_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01555_));
 sky130_fd_sc_hd__o211a_2 _20309_ (.A1(_01553_),
    .A2(_01550_),
    .B1(_09690_),
    .C1(_01555_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00400_));
 sky130_fd_sc_hd__a41oi_2 _20310_ (.A1(\a_l[14] ),
    .A2(\b_l[14] ),
    .A3(\a_l[15] ),
    .A4(\b_l[15] ),
    .B1(_01546_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_01556_));
 sky130_fd_sc_hd__a21oi_2 _20311_ (.A1(_01555_),
    .A2(_01556_),
    .B1(rst),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_00401_));
 sky130_fd_sc_hd__and2_2 _20312_ (.A(_09690_),
    .B(a[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00402_));
 sky130_fd_sc_hd__and2_2 _20313_ (.A(_09690_),
    .B(a[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00403_));
 sky130_fd_sc_hd__and2_2 _20314_ (.A(_09690_),
    .B(a[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00404_));
 sky130_fd_sc_hd__and2_2 _20315_ (.A(_09690_),
    .B(a[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00405_));
 sky130_fd_sc_hd__and2_2 _20316_ (.A(_09690_),
    .B(a[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00406_));
 sky130_fd_sc_hd__and2_2 _20317_ (.A(_09690_),
    .B(a[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00407_));
 sky130_fd_sc_hd__and2_2 _20318_ (.A(_09690_),
    .B(a[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00408_));
 sky130_fd_sc_hd__and2_2 _20319_ (.A(_09690_),
    .B(a[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00409_));
 sky130_fd_sc_hd__and2_2 _20320_ (.A(_09690_),
    .B(a[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00410_));
 sky130_fd_sc_hd__and2_2 _20321_ (.A(_09690_),
    .B(a[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00411_));
 sky130_fd_sc_hd__and2_2 _20322_ (.A(_09690_),
    .B(a[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00412_));
 sky130_fd_sc_hd__and2_2 _20323_ (.A(_09690_),
    .B(a[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00413_));
 sky130_fd_sc_hd__and2_2 _20324_ (.A(_09690_),
    .B(a[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00414_));
 sky130_fd_sc_hd__and2_2 _20325_ (.A(_09690_),
    .B(a[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00415_));
 sky130_fd_sc_hd__and2_2 _20326_ (.A(_09690_),
    .B(a[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00416_));
 sky130_fd_sc_hd__and2_2 _20327_ (.A(_09690_),
    .B(a[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00417_));
 sky130_fd_sc_hd__and2_2 _20328_ (.A(_09690_),
    .B(a[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00418_));
 sky130_fd_sc_hd__and2_2 _20329_ (.A(_09690_),
    .B(a[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00419_));
 sky130_fd_sc_hd__and2_2 _20330_ (.A(_09690_),
    .B(a[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00420_));
 sky130_fd_sc_hd__and2_2 _20331_ (.A(_09690_),
    .B(a[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00421_));
 sky130_fd_sc_hd__and2_2 _20332_ (.A(_09690_),
    .B(a[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00422_));
 sky130_fd_sc_hd__and2_2 _20333_ (.A(_09690_),
    .B(a[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00423_));
 sky130_fd_sc_hd__and2_2 _20334_ (.A(_09690_),
    .B(a[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00424_));
 sky130_fd_sc_hd__and2_2 _20335_ (.A(_09690_),
    .B(a[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00425_));
 sky130_fd_sc_hd__and2_2 _20336_ (.A(_09690_),
    .B(a[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00426_));
 sky130_fd_sc_hd__and2_2 _20337_ (.A(_09690_),
    .B(a[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00427_));
 sky130_fd_sc_hd__and2_2 _20338_ (.A(_09690_),
    .B(a[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00428_));
 sky130_fd_sc_hd__and2_2 _20339_ (.A(_09690_),
    .B(a[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00429_));
 sky130_fd_sc_hd__and2_2 _20340_ (.A(_09690_),
    .B(a[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00430_));
 sky130_fd_sc_hd__and2_2 _20341_ (.A(_09690_),
    .B(a[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00431_));
 sky130_fd_sc_hd__and2_2 _20342_ (.A(_09690_),
    .B(a[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00432_));
 sky130_fd_sc_hd__and2_2 _20343_ (.A(_09690_),
    .B(a[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00433_));
 sky130_fd_sc_hd__and2_2 _20344_ (.A(_09690_),
    .B(b[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00434_));
 sky130_fd_sc_hd__and2_2 _20345_ (.A(_09690_),
    .B(b[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00435_));
 sky130_fd_sc_hd__and2_2 _20346_ (.A(_09690_),
    .B(b[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00436_));
 sky130_fd_sc_hd__and2_2 _20347_ (.A(_09690_),
    .B(b[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00437_));
 sky130_fd_sc_hd__and2_2 _20348_ (.A(_09690_),
    .B(b[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00438_));
 sky130_fd_sc_hd__and2_2 _20349_ (.A(_09690_),
    .B(b[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00439_));
 sky130_fd_sc_hd__and2_2 _20350_ (.A(_09690_),
    .B(b[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00440_));
 sky130_fd_sc_hd__and2_2 _20351_ (.A(_09690_),
    .B(b[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00441_));
 sky130_fd_sc_hd__and2_2 _20352_ (.A(_09690_),
    .B(b[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00442_));
 sky130_fd_sc_hd__and2_2 _20353_ (.A(_09690_),
    .B(b[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00443_));
 sky130_fd_sc_hd__and2_2 _20354_ (.A(_09690_),
    .B(b[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00444_));
 sky130_fd_sc_hd__and2_2 _20355_ (.A(_09690_),
    .B(b[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00445_));
 sky130_fd_sc_hd__and2_2 _20356_ (.A(_09690_),
    .B(b[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00446_));
 sky130_fd_sc_hd__and2_2 _20357_ (.A(_09690_),
    .B(b[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00447_));
 sky130_fd_sc_hd__and2_2 _20358_ (.A(_09690_),
    .B(b[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00448_));
 sky130_fd_sc_hd__and2_2 _20359_ (.A(_09690_),
    .B(b[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_00449_));
 sky130_fd_sc_hd__dfxtp_2 _20360_ (.CLK(clk),
    .D(_00000_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20361_ (.CLK(clk),
    .D(_00001_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20362_ (.CLK(clk),
    .D(_00002_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20363_ (.CLK(clk),
    .D(_00003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20364_ (.CLK(clk),
    .D(_00004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20365_ (.CLK(clk),
    .D(_00005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20366_ (.CLK(clk),
    .D(_00006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20367_ (.CLK(clk),
    .D(_00007_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20368_ (.CLK(clk),
    .D(_00008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20369_ (.CLK(clk),
    .D(_00009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20370_ (.CLK(clk),
    .D(_00010_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20371_ (.CLK(clk),
    .D(_00011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20372_ (.CLK(clk),
    .D(_00012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20373_ (.CLK(clk),
    .D(_00013_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20374_ (.CLK(clk),
    .D(_00014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20375_ (.CLK(clk),
    .D(_00015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_l[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20376_ (.CLK(clk),
    .D(_00016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[0]));
 sky130_fd_sc_hd__dfxtp_2 _20377_ (.CLK(clk),
    .D(_00017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[1]));
 sky130_fd_sc_hd__dfxtp_2 _20378_ (.CLK(clk),
    .D(_00018_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[2]));
 sky130_fd_sc_hd__dfxtp_2 _20379_ (.CLK(clk),
    .D(_00019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[3]));
 sky130_fd_sc_hd__dfxtp_2 _20380_ (.CLK(clk),
    .D(_00020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[4]));
 sky130_fd_sc_hd__dfxtp_2 _20381_ (.CLK(clk),
    .D(_00021_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[5]));
 sky130_fd_sc_hd__dfxtp_2 _20382_ (.CLK(clk),
    .D(_00022_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[6]));
 sky130_fd_sc_hd__dfxtp_2 _20383_ (.CLK(clk),
    .D(_00023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[7]));
 sky130_fd_sc_hd__dfxtp_2 _20384_ (.CLK(clk),
    .D(_00024_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[8]));
 sky130_fd_sc_hd__dfxtp_2 _20385_ (.CLK(clk),
    .D(_00025_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[9]));
 sky130_fd_sc_hd__dfxtp_2 _20386_ (.CLK(clk),
    .D(_00026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[10]));
 sky130_fd_sc_hd__dfxtp_2 _20387_ (.CLK(clk),
    .D(_00027_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[11]));
 sky130_fd_sc_hd__dfxtp_2 _20388_ (.CLK(clk),
    .D(_00028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[12]));
 sky130_fd_sc_hd__dfxtp_2 _20389_ (.CLK(clk),
    .D(_00029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[13]));
 sky130_fd_sc_hd__dfxtp_2 _20390_ (.CLK(clk),
    .D(_00030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[14]));
 sky130_fd_sc_hd__dfxtp_2 _20391_ (.CLK(clk),
    .D(_00031_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[15]));
 sky130_fd_sc_hd__dfxtp_2 _20392_ (.CLK(clk),
    .D(_00032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[16]));
 sky130_fd_sc_hd__dfxtp_2 _20393_ (.CLK(clk),
    .D(_00033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[17]));
 sky130_fd_sc_hd__dfxtp_2 _20394_ (.CLK(clk),
    .D(_00034_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[18]));
 sky130_fd_sc_hd__dfxtp_2 _20395_ (.CLK(clk),
    .D(_00035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[19]));
 sky130_fd_sc_hd__dfxtp_2 _20396_ (.CLK(clk),
    .D(_00036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[20]));
 sky130_fd_sc_hd__dfxtp_2 _20397_ (.CLK(clk),
    .D(_00037_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[21]));
 sky130_fd_sc_hd__dfxtp_2 _20398_ (.CLK(clk),
    .D(_00038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[22]));
 sky130_fd_sc_hd__dfxtp_2 _20399_ (.CLK(clk),
    .D(_00039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[23]));
 sky130_fd_sc_hd__dfxtp_2 _20400_ (.CLK(clk),
    .D(_00040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[24]));
 sky130_fd_sc_hd__dfxtp_2 _20401_ (.CLK(clk),
    .D(_00041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[25]));
 sky130_fd_sc_hd__dfxtp_2 _20402_ (.CLK(clk),
    .D(_00042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[26]));
 sky130_fd_sc_hd__dfxtp_2 _20403_ (.CLK(clk),
    .D(_00043_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[27]));
 sky130_fd_sc_hd__dfxtp_2 _20404_ (.CLK(clk),
    .D(_00044_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[28]));
 sky130_fd_sc_hd__dfxtp_2 _20405_ (.CLK(clk),
    .D(_00045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[29]));
 sky130_fd_sc_hd__dfxtp_2 _20406_ (.CLK(clk),
    .D(_00046_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[30]));
 sky130_fd_sc_hd__dfxtp_2 _20407_ (.CLK(clk),
    .D(_00047_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[31]));
 sky130_fd_sc_hd__dfxtp_2 _20408_ (.CLK(clk),
    .D(_00048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[32]));
 sky130_fd_sc_hd__dfxtp_2 _20409_ (.CLK(clk),
    .D(_00049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[33]));
 sky130_fd_sc_hd__dfxtp_2 _20410_ (.CLK(clk),
    .D(_00050_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[34]));
 sky130_fd_sc_hd__dfxtp_2 _20411_ (.CLK(clk),
    .D(_00051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[35]));
 sky130_fd_sc_hd__dfxtp_2 _20412_ (.CLK(clk),
    .D(_00052_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[36]));
 sky130_fd_sc_hd__dfxtp_2 _20413_ (.CLK(clk),
    .D(_00053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[37]));
 sky130_fd_sc_hd__dfxtp_2 _20414_ (.CLK(clk),
    .D(_00054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[38]));
 sky130_fd_sc_hd__dfxtp_2 _20415_ (.CLK(clk),
    .D(_00055_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[39]));
 sky130_fd_sc_hd__dfxtp_2 _20416_ (.CLK(clk),
    .D(_00056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[40]));
 sky130_fd_sc_hd__dfxtp_2 _20417_ (.CLK(clk),
    .D(_00057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[41]));
 sky130_fd_sc_hd__dfxtp_2 _20418_ (.CLK(clk),
    .D(_00058_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[42]));
 sky130_fd_sc_hd__dfxtp_2 _20419_ (.CLK(clk),
    .D(_00059_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[43]));
 sky130_fd_sc_hd__dfxtp_2 _20420_ (.CLK(clk),
    .D(_00060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[44]));
 sky130_fd_sc_hd__dfxtp_2 _20421_ (.CLK(clk),
    .D(_00061_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[45]));
 sky130_fd_sc_hd__dfxtp_2 _20422_ (.CLK(clk),
    .D(_00062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[46]));
 sky130_fd_sc_hd__dfxtp_2 _20423_ (.CLK(clk),
    .D(_00063_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[47]));
 sky130_fd_sc_hd__dfxtp_2 _20424_ (.CLK(clk),
    .D(_00064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[48]));
 sky130_fd_sc_hd__dfxtp_2 _20425_ (.CLK(clk),
    .D(_00065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[49]));
 sky130_fd_sc_hd__dfxtp_2 _20426_ (.CLK(clk),
    .D(_00066_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[50]));
 sky130_fd_sc_hd__dfxtp_2 _20427_ (.CLK(clk),
    .D(_00067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[51]));
 sky130_fd_sc_hd__dfxtp_2 _20428_ (.CLK(clk),
    .D(_00068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[52]));
 sky130_fd_sc_hd__dfxtp_2 _20429_ (.CLK(clk),
    .D(_00069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[53]));
 sky130_fd_sc_hd__dfxtp_2 _20430_ (.CLK(clk),
    .D(_00070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[54]));
 sky130_fd_sc_hd__dfxtp_2 _20431_ (.CLK(clk),
    .D(_00071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[55]));
 sky130_fd_sc_hd__dfxtp_2 _20432_ (.CLK(clk),
    .D(_00072_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[56]));
 sky130_fd_sc_hd__dfxtp_2 _20433_ (.CLK(clk),
    .D(_00073_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[57]));
 sky130_fd_sc_hd__dfxtp_2 _20434_ (.CLK(clk),
    .D(_00074_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[58]));
 sky130_fd_sc_hd__dfxtp_2 _20435_ (.CLK(clk),
    .D(_00075_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[59]));
 sky130_fd_sc_hd__dfxtp_2 _20436_ (.CLK(clk),
    .D(_00076_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[60]));
 sky130_fd_sc_hd__dfxtp_2 _20437_ (.CLK(clk),
    .D(_00077_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[61]));
 sky130_fd_sc_hd__dfxtp_2 _20438_ (.CLK(clk),
    .D(_00078_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[62]));
 sky130_fd_sc_hd__dfxtp_2 _20439_ (.CLK(clk),
    .D(_00079_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(p[63]));
 sky130_fd_sc_hd__dfxtp_2 _20440_ (.CLK(clk),
    .D(_00080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[32] ));
 sky130_fd_sc_hd__dfxtp_2 _20441_ (.CLK(clk),
    .D(_00081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[33] ));
 sky130_fd_sc_hd__dfxtp_2 _20442_ (.CLK(clk),
    .D(_00082_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[34] ));
 sky130_fd_sc_hd__dfxtp_2 _20443_ (.CLK(clk),
    .D(_00083_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[35] ));
 sky130_fd_sc_hd__dfxtp_2 _20444_ (.CLK(clk),
    .D(_00084_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[36] ));
 sky130_fd_sc_hd__dfxtp_2 _20445_ (.CLK(clk),
    .D(_00085_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[37] ));
 sky130_fd_sc_hd__dfxtp_2 _20446_ (.CLK(clk),
    .D(_00086_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[38] ));
 sky130_fd_sc_hd__dfxtp_2 _20447_ (.CLK(clk),
    .D(_00087_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[39] ));
 sky130_fd_sc_hd__dfxtp_2 _20448_ (.CLK(clk),
    .D(_00088_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[40] ));
 sky130_fd_sc_hd__dfxtp_2 _20449_ (.CLK(clk),
    .D(_00089_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[41] ));
 sky130_fd_sc_hd__dfxtp_2 _20450_ (.CLK(clk),
    .D(_00090_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[42] ));
 sky130_fd_sc_hd__dfxtp_2 _20451_ (.CLK(clk),
    .D(_00091_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[43] ));
 sky130_fd_sc_hd__dfxtp_2 _20452_ (.CLK(clk),
    .D(_00092_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[44] ));
 sky130_fd_sc_hd__dfxtp_2 _20453_ (.CLK(clk),
    .D(_00093_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[45] ));
 sky130_fd_sc_hd__dfxtp_2 _20454_ (.CLK(clk),
    .D(_00094_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[46] ));
 sky130_fd_sc_hd__dfxtp_2 _20455_ (.CLK(clk),
    .D(_00095_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[47] ));
 sky130_fd_sc_hd__dfxtp_2 _20456_ (.CLK(clk),
    .D(_00096_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[48] ));
 sky130_fd_sc_hd__dfxtp_2 _20457_ (.CLK(clk),
    .D(_00097_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[49] ));
 sky130_fd_sc_hd__dfxtp_2 _20458_ (.CLK(clk),
    .D(_00098_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[50] ));
 sky130_fd_sc_hd__dfxtp_2 _20459_ (.CLK(clk),
    .D(_00099_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[51] ));
 sky130_fd_sc_hd__dfxtp_2 _20460_ (.CLK(clk),
    .D(_00100_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[52] ));
 sky130_fd_sc_hd__dfxtp_2 _20461_ (.CLK(clk),
    .D(_00101_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[53] ));
 sky130_fd_sc_hd__dfxtp_2 _20462_ (.CLK(clk),
    .D(_00102_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[54] ));
 sky130_fd_sc_hd__dfxtp_2 _20463_ (.CLK(clk),
    .D(_00103_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[55] ));
 sky130_fd_sc_hd__dfxtp_2 _20464_ (.CLK(clk),
    .D(_00104_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[56] ));
 sky130_fd_sc_hd__dfxtp_2 _20465_ (.CLK(clk),
    .D(_00105_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[57] ));
 sky130_fd_sc_hd__dfxtp_2 _20466_ (.CLK(clk),
    .D(_00106_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[58] ));
 sky130_fd_sc_hd__dfxtp_2 _20467_ (.CLK(clk),
    .D(_00107_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[59] ));
 sky130_fd_sc_hd__dfxtp_2 _20468_ (.CLK(clk),
    .D(_00108_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[60] ));
 sky130_fd_sc_hd__dfxtp_2 _20469_ (.CLK(clk),
    .D(_00109_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[61] ));
 sky130_fd_sc_hd__dfxtp_2 _20470_ (.CLK(clk),
    .D(_00110_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[62] ));
 sky130_fd_sc_hd__dfxtp_2 _20471_ (.CLK(clk),
    .D(_00111_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_high[63] ));
 sky130_fd_sc_hd__dfxtp_2 _20472_ (.CLK(clk),
    .D(_00112_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20473_ (.CLK(clk),
    .D(_00113_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20474_ (.CLK(clk),
    .D(_00114_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20475_ (.CLK(clk),
    .D(_00115_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20476_ (.CLK(clk),
    .D(_00116_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20477_ (.CLK(clk),
    .D(_00117_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20478_ (.CLK(clk),
    .D(_00118_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20479_ (.CLK(clk),
    .D(_00119_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20480_ (.CLK(clk),
    .D(_00120_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20481_ (.CLK(clk),
    .D(_00121_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20482_ (.CLK(clk),
    .D(_00122_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20483_ (.CLK(clk),
    .D(_00123_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20484_ (.CLK(clk),
    .D(_00124_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20485_ (.CLK(clk),
    .D(_00125_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20486_ (.CLK(clk),
    .D(_00126_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20487_ (.CLK(clk),
    .D(_00127_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20488_ (.CLK(clk),
    .D(_00128_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[32] ));
 sky130_fd_sc_hd__dfxtp_2 _20489_ (.CLK(clk),
    .D(_00129_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[33] ));
 sky130_fd_sc_hd__dfxtp_2 _20490_ (.CLK(clk),
    .D(_00130_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[34] ));
 sky130_fd_sc_hd__dfxtp_2 _20491_ (.CLK(clk),
    .D(_00131_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[35] ));
 sky130_fd_sc_hd__dfxtp_2 _20492_ (.CLK(clk),
    .D(_00132_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[36] ));
 sky130_fd_sc_hd__dfxtp_2 _20493_ (.CLK(clk),
    .D(_00133_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[37] ));
 sky130_fd_sc_hd__dfxtp_2 _20494_ (.CLK(clk),
    .D(_00134_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[38] ));
 sky130_fd_sc_hd__dfxtp_2 _20495_ (.CLK(clk),
    .D(_00135_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[39] ));
 sky130_fd_sc_hd__dfxtp_2 _20496_ (.CLK(clk),
    .D(_00136_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[40] ));
 sky130_fd_sc_hd__dfxtp_2 _20497_ (.CLK(clk),
    .D(_00137_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[41] ));
 sky130_fd_sc_hd__dfxtp_2 _20498_ (.CLK(clk),
    .D(_00138_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[42] ));
 sky130_fd_sc_hd__dfxtp_2 _20499_ (.CLK(clk),
    .D(_00139_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[43] ));
 sky130_fd_sc_hd__dfxtp_2 _20500_ (.CLK(clk),
    .D(_00140_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[44] ));
 sky130_fd_sc_hd__dfxtp_2 _20501_ (.CLK(clk),
    .D(_00141_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[45] ));
 sky130_fd_sc_hd__dfxtp_2 _20502_ (.CLK(clk),
    .D(_00142_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[46] ));
 sky130_fd_sc_hd__dfxtp_2 _20503_ (.CLK(clk),
    .D(_00143_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[47] ));
 sky130_fd_sc_hd__dfxtp_2 _20504_ (.CLK(clk),
    .D(_00144_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_mid[48] ));
 sky130_fd_sc_hd__dfxtp_2 _20505_ (.CLK(clk),
    .D(_00145_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20506_ (.CLK(clk),
    .D(_00146_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20507_ (.CLK(clk),
    .D(_00147_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20508_ (.CLK(clk),
    .D(_00148_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20509_ (.CLK(clk),
    .D(_00149_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20510_ (.CLK(clk),
    .D(_00150_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20511_ (.CLK(clk),
    .D(_00151_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20512_ (.CLK(clk),
    .D(_00152_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20513_ (.CLK(clk),
    .D(_00153_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20514_ (.CLK(clk),
    .D(_00154_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20515_ (.CLK(clk),
    .D(_00155_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20516_ (.CLK(clk),
    .D(_00156_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20517_ (.CLK(clk),
    .D(_00157_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20518_ (.CLK(clk),
    .D(_00158_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20519_ (.CLK(clk),
    .D(_00159_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20520_ (.CLK(clk),
    .D(_00160_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20521_ (.CLK(clk),
    .D(_00161_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20522_ (.CLK(clk),
    .D(_00162_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20523_ (.CLK(clk),
    .D(_00163_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20524_ (.CLK(clk),
    .D(_00164_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20525_ (.CLK(clk),
    .D(_00165_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20526_ (.CLK(clk),
    .D(_00166_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20527_ (.CLK(clk),
    .D(_00167_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20528_ (.CLK(clk),
    .D(_00168_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20529_ (.CLK(clk),
    .D(_00169_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20530_ (.CLK(clk),
    .D(_00170_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20531_ (.CLK(clk),
    .D(_00171_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20532_ (.CLK(clk),
    .D(_00172_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20533_ (.CLK(clk),
    .D(_00173_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20534_ (.CLK(clk),
    .D(_00174_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20535_ (.CLK(clk),
    .D(_00175_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20536_ (.CLK(clk),
    .D(_00176_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\term_low[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20537_ (.CLK(clk),
    .D(_00177_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20538_ (.CLK(clk),
    .D(_00178_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20539_ (.CLK(clk),
    .D(_00179_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20540_ (.CLK(clk),
    .D(_00180_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20541_ (.CLK(clk),
    .D(_00181_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20542_ (.CLK(clk),
    .D(_00182_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20543_ (.CLK(clk),
    .D(_00183_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20544_ (.CLK(clk),
    .D(_00184_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20545_ (.CLK(clk),
    .D(_00185_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20546_ (.CLK(clk),
    .D(_00186_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20547_ (.CLK(clk),
    .D(_00187_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20548_ (.CLK(clk),
    .D(_00188_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20549_ (.CLK(clk),
    .D(_00189_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20550_ (.CLK(clk),
    .D(_00190_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20551_ (.CLK(clk),
    .D(_00191_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20552_ (.CLK(clk),
    .D(_00192_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20553_ (.CLK(clk),
    .D(_00193_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20554_ (.CLK(clk),
    .D(_00194_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20555_ (.CLK(clk),
    .D(_00195_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20556_ (.CLK(clk),
    .D(_00196_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20557_ (.CLK(clk),
    .D(_00197_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20558_ (.CLK(clk),
    .D(_00198_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20559_ (.CLK(clk),
    .D(_00199_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20560_ (.CLK(clk),
    .D(_00200_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20561_ (.CLK(clk),
    .D(_00201_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20562_ (.CLK(clk),
    .D(_00202_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20563_ (.CLK(clk),
    .D(_00203_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20564_ (.CLK(clk),
    .D(_00204_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20565_ (.CLK(clk),
    .D(_00205_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20566_ (.CLK(clk),
    .D(_00206_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20567_ (.CLK(clk),
    .D(_00207_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20568_ (.CLK(clk),
    .D(_00208_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20569_ (.CLK(clk),
    .D(_00209_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\mid_sum[32] ));
 sky130_fd_sc_hd__dfxtp_2 _20570_ (.CLK(clk),
    .D(_00210_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20571_ (.CLK(clk),
    .D(_00211_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20572_ (.CLK(clk),
    .D(_00212_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20573_ (.CLK(clk),
    .D(_00213_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20574_ (.CLK(clk),
    .D(_00214_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20575_ (.CLK(clk),
    .D(_00215_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20576_ (.CLK(clk),
    .D(_00216_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20577_ (.CLK(clk),
    .D(_00217_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20578_ (.CLK(clk),
    .D(_00218_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20579_ (.CLK(clk),
    .D(_00219_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20580_ (.CLK(clk),
    .D(_00220_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20581_ (.CLK(clk),
    .D(_00221_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20582_ (.CLK(clk),
    .D(_00222_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20583_ (.CLK(clk),
    .D(_00223_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20584_ (.CLK(clk),
    .D(_00224_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20585_ (.CLK(clk),
    .D(_00225_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20586_ (.CLK(clk),
    .D(_00226_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20587_ (.CLK(clk),
    .D(_00227_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20588_ (.CLK(clk),
    .D(_00228_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20589_ (.CLK(clk),
    .D(_00229_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20590_ (.CLK(clk),
    .D(_00230_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20591_ (.CLK(clk),
    .D(_00231_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20592_ (.CLK(clk),
    .D(_00232_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20593_ (.CLK(clk),
    .D(_00233_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20594_ (.CLK(clk),
    .D(_00234_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20595_ (.CLK(clk),
    .D(_00235_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20596_ (.CLK(clk),
    .D(_00236_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20597_ (.CLK(clk),
    .D(_00237_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20598_ (.CLK(clk),
    .D(_00238_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20599_ (.CLK(clk),
    .D(_00239_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20600_ (.CLK(clk),
    .D(_00240_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20601_ (.CLK(clk),
    .D(_00241_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh_pipe[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20602_ (.CLK(clk),
    .D(_00242_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20603_ (.CLK(clk),
    .D(_00243_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20604_ (.CLK(clk),
    .D(_00244_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20605_ (.CLK(clk),
    .D(_00245_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20606_ (.CLK(clk),
    .D(_00246_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20607_ (.CLK(clk),
    .D(_00247_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20608_ (.CLK(clk),
    .D(_00248_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20609_ (.CLK(clk),
    .D(_00249_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20610_ (.CLK(clk),
    .D(_00250_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20611_ (.CLK(clk),
    .D(_00251_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20612_ (.CLK(clk),
    .D(_00252_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20613_ (.CLK(clk),
    .D(_00253_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20614_ (.CLK(clk),
    .D(_00254_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20615_ (.CLK(clk),
    .D(_00255_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20616_ (.CLK(clk),
    .D(_00256_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20617_ (.CLK(clk),
    .D(_00257_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20618_ (.CLK(clk),
    .D(_00258_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20619_ (.CLK(clk),
    .D(_00259_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20620_ (.CLK(clk),
    .D(_00260_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20621_ (.CLK(clk),
    .D(_00261_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20622_ (.CLK(clk),
    .D(_00262_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20623_ (.CLK(clk),
    .D(_00263_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20624_ (.CLK(clk),
    .D(_00264_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20625_ (.CLK(clk),
    .D(_00265_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20626_ (.CLK(clk),
    .D(_00266_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20627_ (.CLK(clk),
    .D(_00267_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20628_ (.CLK(clk),
    .D(_00268_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20629_ (.CLK(clk),
    .D(_00269_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20630_ (.CLK(clk),
    .D(_00270_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20631_ (.CLK(clk),
    .D(_00271_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20632_ (.CLK(clk),
    .D(_00272_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20633_ (.CLK(clk),
    .D(_00273_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll_pipe[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20634_ (.CLK(clk),
    .D(_00274_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20635_ (.CLK(clk),
    .D(_00275_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20636_ (.CLK(clk),
    .D(_00276_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20637_ (.CLK(clk),
    .D(_00277_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20638_ (.CLK(clk),
    .D(_00278_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20639_ (.CLK(clk),
    .D(_00279_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20640_ (.CLK(clk),
    .D(_00280_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20641_ (.CLK(clk),
    .D(_00281_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20642_ (.CLK(clk),
    .D(_00282_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20643_ (.CLK(clk),
    .D(_00283_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20644_ (.CLK(clk),
    .D(_00284_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20645_ (.CLK(clk),
    .D(_00285_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20646_ (.CLK(clk),
    .D(_00286_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20647_ (.CLK(clk),
    .D(_00287_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20648_ (.CLK(clk),
    .D(_00288_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20649_ (.CLK(clk),
    .D(_00289_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20650_ (.CLK(clk),
    .D(_00290_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20651_ (.CLK(clk),
    .D(_00291_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20652_ (.CLK(clk),
    .D(_00292_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20653_ (.CLK(clk),
    .D(_00293_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20654_ (.CLK(clk),
    .D(_00294_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20655_ (.CLK(clk),
    .D(_00295_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20656_ (.CLK(clk),
    .D(_00296_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20657_ (.CLK(clk),
    .D(_00297_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20658_ (.CLK(clk),
    .D(_00298_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20659_ (.CLK(clk),
    .D(_00299_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20660_ (.CLK(clk),
    .D(_00300_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20661_ (.CLK(clk),
    .D(_00301_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20662_ (.CLK(clk),
    .D(_00302_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20663_ (.CLK(clk),
    .D(_00303_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20664_ (.CLK(clk),
    .D(_00304_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20665_ (.CLK(clk),
    .D(_00305_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hh[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20666_ (.CLK(clk),
    .D(_00306_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20667_ (.CLK(clk),
    .D(_00307_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20668_ (.CLK(clk),
    .D(_00308_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20669_ (.CLK(clk),
    .D(_00309_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20670_ (.CLK(clk),
    .D(_00310_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20671_ (.CLK(clk),
    .D(_00311_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20672_ (.CLK(clk),
    .D(_00312_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20673_ (.CLK(clk),
    .D(_00313_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20674_ (.CLK(clk),
    .D(_00314_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20675_ (.CLK(clk),
    .D(_00315_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20676_ (.CLK(clk),
    .D(_00316_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20677_ (.CLK(clk),
    .D(_00317_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20678_ (.CLK(clk),
    .D(_00318_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20679_ (.CLK(clk),
    .D(_00319_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20680_ (.CLK(clk),
    .D(_00320_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20681_ (.CLK(clk),
    .D(_00321_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20682_ (.CLK(clk),
    .D(_00322_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20683_ (.CLK(clk),
    .D(_00323_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20684_ (.CLK(clk),
    .D(_00324_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20685_ (.CLK(clk),
    .D(_00325_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20686_ (.CLK(clk),
    .D(_00326_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20687_ (.CLK(clk),
    .D(_00327_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20688_ (.CLK(clk),
    .D(_00328_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20689_ (.CLK(clk),
    .D(_00329_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20690_ (.CLK(clk),
    .D(_00330_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20691_ (.CLK(clk),
    .D(_00331_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20692_ (.CLK(clk),
    .D(_00332_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20693_ (.CLK(clk),
    .D(_00333_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20694_ (.CLK(clk),
    .D(_00334_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20695_ (.CLK(clk),
    .D(_00335_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20696_ (.CLK(clk),
    .D(_00336_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20697_ (.CLK(clk),
    .D(_00337_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_hl[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20698_ (.CLK(clk),
    .D(_00338_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20699_ (.CLK(clk),
    .D(_00339_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20700_ (.CLK(clk),
    .D(_00340_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20701_ (.CLK(clk),
    .D(_00341_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20702_ (.CLK(clk),
    .D(_00342_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20703_ (.CLK(clk),
    .D(_00343_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20704_ (.CLK(clk),
    .D(_00344_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20705_ (.CLK(clk),
    .D(_00345_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20706_ (.CLK(clk),
    .D(_00346_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20707_ (.CLK(clk),
    .D(_00347_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20708_ (.CLK(clk),
    .D(_00348_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20709_ (.CLK(clk),
    .D(_00349_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20710_ (.CLK(clk),
    .D(_00350_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20711_ (.CLK(clk),
    .D(_00351_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20712_ (.CLK(clk),
    .D(_00352_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20713_ (.CLK(clk),
    .D(_00353_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20714_ (.CLK(clk),
    .D(_00354_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20715_ (.CLK(clk),
    .D(_00355_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20716_ (.CLK(clk),
    .D(_00356_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20717_ (.CLK(clk),
    .D(_00357_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20718_ (.CLK(clk),
    .D(_00358_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20719_ (.CLK(clk),
    .D(_00359_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20720_ (.CLK(clk),
    .D(_00360_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20721_ (.CLK(clk),
    .D(_00361_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20722_ (.CLK(clk),
    .D(_00362_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20723_ (.CLK(clk),
    .D(_00363_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20724_ (.CLK(clk),
    .D(_00364_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20725_ (.CLK(clk),
    .D(_00365_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20726_ (.CLK(clk),
    .D(_00366_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20727_ (.CLK(clk),
    .D(_00367_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20728_ (.CLK(clk),
    .D(_00368_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20729_ (.CLK(clk),
    .D(_00369_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_lh[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20730_ (.CLK(clk),
    .D(_00370_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20731_ (.CLK(clk),
    .D(_00371_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20732_ (.CLK(clk),
    .D(_00372_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20733_ (.CLK(clk),
    .D(_00373_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20734_ (.CLK(clk),
    .D(_00374_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20735_ (.CLK(clk),
    .D(_00375_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20736_ (.CLK(clk),
    .D(_00376_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20737_ (.CLK(clk),
    .D(_00377_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20738_ (.CLK(clk),
    .D(_00378_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20739_ (.CLK(clk),
    .D(_00379_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20740_ (.CLK(clk),
    .D(_00380_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20741_ (.CLK(clk),
    .D(_00381_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20742_ (.CLK(clk),
    .D(_00382_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20743_ (.CLK(clk),
    .D(_00383_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20744_ (.CLK(clk),
    .D(_00384_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20745_ (.CLK(clk),
    .D(_00385_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20746_ (.CLK(clk),
    .D(_00386_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[16] ));
 sky130_fd_sc_hd__dfxtp_2 _20747_ (.CLK(clk),
    .D(_00387_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[17] ));
 sky130_fd_sc_hd__dfxtp_2 _20748_ (.CLK(clk),
    .D(_00388_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[18] ));
 sky130_fd_sc_hd__dfxtp_2 _20749_ (.CLK(clk),
    .D(_00389_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[19] ));
 sky130_fd_sc_hd__dfxtp_2 _20750_ (.CLK(clk),
    .D(_00390_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[20] ));
 sky130_fd_sc_hd__dfxtp_2 _20751_ (.CLK(clk),
    .D(_00391_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[21] ));
 sky130_fd_sc_hd__dfxtp_2 _20752_ (.CLK(clk),
    .D(_00392_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[22] ));
 sky130_fd_sc_hd__dfxtp_2 _20753_ (.CLK(clk),
    .D(_00393_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[23] ));
 sky130_fd_sc_hd__dfxtp_2 _20754_ (.CLK(clk),
    .D(_00394_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[24] ));
 sky130_fd_sc_hd__dfxtp_2 _20755_ (.CLK(clk),
    .D(_00395_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[25] ));
 sky130_fd_sc_hd__dfxtp_2 _20756_ (.CLK(clk),
    .D(_00396_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[26] ));
 sky130_fd_sc_hd__dfxtp_2 _20757_ (.CLK(clk),
    .D(_00397_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[27] ));
 sky130_fd_sc_hd__dfxtp_2 _20758_ (.CLK(clk),
    .D(_00398_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[28] ));
 sky130_fd_sc_hd__dfxtp_2 _20759_ (.CLK(clk),
    .D(_00399_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[29] ));
 sky130_fd_sc_hd__dfxtp_2 _20760_ (.CLK(clk),
    .D(_00400_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[30] ));
 sky130_fd_sc_hd__dfxtp_2 _20761_ (.CLK(clk),
    .D(_00401_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\p_ll[31] ));
 sky130_fd_sc_hd__dfxtp_2 _20762_ (.CLK(clk),
    .D(_00402_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20763_ (.CLK(clk),
    .D(_00403_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20764_ (.CLK(clk),
    .D(_00404_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20765_ (.CLK(clk),
    .D(_00405_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20766_ (.CLK(clk),
    .D(_00406_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20767_ (.CLK(clk),
    .D(_00407_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20768_ (.CLK(clk),
    .D(_00408_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20769_ (.CLK(clk),
    .D(_00409_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20770_ (.CLK(clk),
    .D(_00410_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20771_ (.CLK(clk),
    .D(_00411_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20772_ (.CLK(clk),
    .D(_00412_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20773_ (.CLK(clk),
    .D(_00413_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20774_ (.CLK(clk),
    .D(_00414_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20775_ (.CLK(clk),
    .D(_00415_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20776_ (.CLK(clk),
    .D(_00416_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20777_ (.CLK(clk),
    .D(_00417_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_h[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20778_ (.CLK(clk),
    .D(_00418_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20779_ (.CLK(clk),
    .D(_00419_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20780_ (.CLK(clk),
    .D(_00420_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20781_ (.CLK(clk),
    .D(_00421_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20782_ (.CLK(clk),
    .D(_00422_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20783_ (.CLK(clk),
    .D(_00423_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20784_ (.CLK(clk),
    .D(_00424_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20785_ (.CLK(clk),
    .D(_00425_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20786_ (.CLK(clk),
    .D(_00426_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20787_ (.CLK(clk),
    .D(_00427_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20788_ (.CLK(clk),
    .D(_00428_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20789_ (.CLK(clk),
    .D(_00429_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20790_ (.CLK(clk),
    .D(_00430_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20791_ (.CLK(clk),
    .D(_00431_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20792_ (.CLK(clk),
    .D(_00432_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20793_ (.CLK(clk),
    .D(_00433_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\a_l[15] ));
 sky130_fd_sc_hd__dfxtp_2 _20794_ (.CLK(clk),
    .D(_00434_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[0] ));
 sky130_fd_sc_hd__dfxtp_2 _20795_ (.CLK(clk),
    .D(_00435_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[1] ));
 sky130_fd_sc_hd__dfxtp_2 _20796_ (.CLK(clk),
    .D(_00436_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[2] ));
 sky130_fd_sc_hd__dfxtp_2 _20797_ (.CLK(clk),
    .D(_00437_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[3] ));
 sky130_fd_sc_hd__dfxtp_2 _20798_ (.CLK(clk),
    .D(_00438_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[4] ));
 sky130_fd_sc_hd__dfxtp_2 _20799_ (.CLK(clk),
    .D(_00439_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[5] ));
 sky130_fd_sc_hd__dfxtp_2 _20800_ (.CLK(clk),
    .D(_00440_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[6] ));
 sky130_fd_sc_hd__dfxtp_2 _20801_ (.CLK(clk),
    .D(_00441_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[7] ));
 sky130_fd_sc_hd__dfxtp_2 _20802_ (.CLK(clk),
    .D(_00442_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[8] ));
 sky130_fd_sc_hd__dfxtp_2 _20803_ (.CLK(clk),
    .D(_00443_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[9] ));
 sky130_fd_sc_hd__dfxtp_2 _20804_ (.CLK(clk),
    .D(_00444_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[10] ));
 sky130_fd_sc_hd__dfxtp_2 _20805_ (.CLK(clk),
    .D(_00445_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[11] ));
 sky130_fd_sc_hd__dfxtp_2 _20806_ (.CLK(clk),
    .D(_00446_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[12] ));
 sky130_fd_sc_hd__dfxtp_2 _20807_ (.CLK(clk),
    .D(_00447_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[13] ));
 sky130_fd_sc_hd__dfxtp_2 _20808_ (.CLK(clk),
    .D(_00448_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[14] ));
 sky130_fd_sc_hd__dfxtp_2 _20809_ (.CLK(clk),
    .D(_00449_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\b_h[15] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_282 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_3010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_3033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_3055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_4000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_4023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_4045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_4068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_5013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5238 (.VGND(VGND),
    .VPWR(VPWR));
endmodule
