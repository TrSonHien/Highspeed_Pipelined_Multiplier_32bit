VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.340 10.640 75.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.340 10.640 125.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.340 10.640 175.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.340 10.640 225.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.340 10.640 275.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.340 10.640 325.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.340 10.640 425.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.340 10.640 475.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.340 10.640 525.940 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.340 10.640 575.940 587.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 594.560 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.030 594.560 81.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 130.030 594.560 131.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 180.030 594.560 181.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 230.030 594.560 231.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 280.030 594.560 281.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 330.030 594.560 331.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 594.560 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 430.030 594.560 431.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 480.030 594.560 481.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 530.030 594.560 531.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 580.030 594.560 581.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 587.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 594.560 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.730 594.560 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 126.730 594.560 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 176.730 594.560 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 226.730 594.560 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 276.730 594.560 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 326.730 594.560 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 594.560 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 426.730 594.560 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 476.730 594.560 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 526.730 594.560 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 576.730 594.560 578.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 413.480 600.000 414.080 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 236.680 600.000 237.280 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 254.360 600.000 254.960 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 272.040 600.000 272.640 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 289.720 600.000 290.320 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 307.400 600.000 308.000 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 325.080 600.000 325.680 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 342.760 600.000 343.360 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 360.440 600.000 361.040 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 378.120 600.000 378.720 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 395.800 600.000 396.400 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 431.160 600.000 431.760 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 59.880 600.000 60.480 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 77.560 600.000 78.160 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 95.240 600.000 95.840 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 112.920 600.000 113.520 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 130.600 600.000 131.200 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 148.280 600.000 148.880 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 165.960 600.000 166.560 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 183.640 600.000 184.240 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 201.320 600.000 201.920 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 219.000 600.000 219.600 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 448.840 600.000 449.440 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 24.520 600.000 25.120 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 42.200 600.000 42.800 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 455.950 596.000 456.230 600.000 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 474.350 596.000 474.630 600.000 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 492.750 596.000 493.030 600.000 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 511.150 596.000 511.430 600.000 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 529.550 596.000 529.830 600.000 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 547.950 596.000 548.230 600.000 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 566.350 596.000 566.630 600.000 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 584.750 596.000 585.030 600.000 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 466.520 600.000 467.120 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 271.950 596.000 272.230 600.000 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 290.350 596.000 290.630 600.000 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 308.750 596.000 309.030 600.000 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 327.150 596.000 327.430 600.000 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 345.550 596.000 345.830 600.000 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 363.950 596.000 364.230 600.000 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 382.350 596.000 382.630 600.000 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 400.750 596.000 401.030 600.000 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 419.150 596.000 419.430 600.000 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 437.550 596.000 437.830 600.000 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 484.200 600.000 484.800 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.950 596.000 88.230 600.000 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 596.000 106.630 600.000 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.750 596.000 125.030 600.000 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.150 596.000 143.430 600.000 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.550 596.000 161.830 600.000 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.950 596.000 180.230 600.000 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 596.000 198.630 600.000 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 216.750 596.000 217.030 600.000 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 596.000 235.430 600.000 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 253.550 596.000 253.830 600.000 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 501.880 600.000 502.480 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 14.350 596.000 14.630 600.000 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 596.000 33.030 600.000 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.150 596.000 51.430 600.000 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.550 596.000 69.830 600.000 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 519.560 600.000 520.160 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 537.240 600.000 537.840 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 554.920 600.000 555.520 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 572.600 600.000 573.200 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 594.510 587.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 4.210 10.640 594.620 587.760 ;
      LAYER met2 ;
        RECT 4.230 595.720 14.070 596.770 ;
        RECT 14.910 595.720 32.470 596.770 ;
        RECT 33.310 595.720 50.870 596.770 ;
        RECT 51.710 595.720 69.270 596.770 ;
        RECT 70.110 595.720 87.670 596.770 ;
        RECT 88.510 595.720 106.070 596.770 ;
        RECT 106.910 595.720 124.470 596.770 ;
        RECT 125.310 595.720 142.870 596.770 ;
        RECT 143.710 595.720 161.270 596.770 ;
        RECT 162.110 595.720 179.670 596.770 ;
        RECT 180.510 595.720 198.070 596.770 ;
        RECT 198.910 595.720 216.470 596.770 ;
        RECT 217.310 595.720 234.870 596.770 ;
        RECT 235.710 595.720 253.270 596.770 ;
        RECT 254.110 595.720 271.670 596.770 ;
        RECT 272.510 595.720 290.070 596.770 ;
        RECT 290.910 595.720 308.470 596.770 ;
        RECT 309.310 595.720 326.870 596.770 ;
        RECT 327.710 595.720 345.270 596.770 ;
        RECT 346.110 595.720 363.670 596.770 ;
        RECT 364.510 595.720 382.070 596.770 ;
        RECT 382.910 595.720 400.470 596.770 ;
        RECT 401.310 595.720 418.870 596.770 ;
        RECT 419.710 595.720 437.270 596.770 ;
        RECT 438.110 595.720 455.670 596.770 ;
        RECT 456.510 595.720 474.070 596.770 ;
        RECT 474.910 595.720 492.470 596.770 ;
        RECT 493.310 595.720 510.870 596.770 ;
        RECT 511.710 595.720 529.270 596.770 ;
        RECT 530.110 595.720 547.670 596.770 ;
        RECT 548.510 595.720 566.070 596.770 ;
        RECT 566.910 595.720 584.470 596.770 ;
        RECT 585.310 595.720 593.760 596.770 ;
        RECT 4.230 4.280 593.760 595.720 ;
        RECT 4.230 4.000 12.230 4.280 ;
        RECT 13.070 4.000 30.170 4.280 ;
        RECT 31.010 4.000 48.110 4.280 ;
        RECT 48.950 4.000 66.050 4.280 ;
        RECT 66.890 4.000 83.990 4.280 ;
        RECT 84.830 4.000 101.930 4.280 ;
        RECT 102.770 4.000 119.870 4.280 ;
        RECT 120.710 4.000 137.810 4.280 ;
        RECT 138.650 4.000 155.750 4.280 ;
        RECT 156.590 4.000 173.690 4.280 ;
        RECT 174.530 4.000 191.630 4.280 ;
        RECT 192.470 4.000 209.570 4.280 ;
        RECT 210.410 4.000 227.510 4.280 ;
        RECT 228.350 4.000 245.450 4.280 ;
        RECT 246.290 4.000 263.390 4.280 ;
        RECT 264.230 4.000 281.330 4.280 ;
        RECT 282.170 4.000 299.270 4.280 ;
        RECT 300.110 4.000 317.210 4.280 ;
        RECT 318.050 4.000 335.150 4.280 ;
        RECT 335.990 4.000 353.090 4.280 ;
        RECT 353.930 4.000 371.030 4.280 ;
        RECT 371.870 4.000 388.970 4.280 ;
        RECT 389.810 4.000 406.910 4.280 ;
        RECT 407.750 4.000 424.850 4.280 ;
        RECT 425.690 4.000 442.790 4.280 ;
        RECT 443.630 4.000 460.730 4.280 ;
        RECT 461.570 4.000 478.670 4.280 ;
        RECT 479.510 4.000 496.610 4.280 ;
        RECT 497.450 4.000 514.550 4.280 ;
        RECT 515.390 4.000 532.490 4.280 ;
        RECT 533.330 4.000 550.430 4.280 ;
        RECT 551.270 4.000 568.370 4.280 ;
        RECT 569.210 4.000 586.310 4.280 ;
        RECT 587.150 4.000 593.760 4.280 ;
      LAYER met3 ;
        RECT 3.990 583.120 596.000 587.685 ;
        RECT 4.400 581.720 596.000 583.120 ;
        RECT 3.990 573.600 596.000 581.720 ;
        RECT 3.990 572.200 595.600 573.600 ;
        RECT 3.990 565.440 596.000 572.200 ;
        RECT 4.400 564.040 596.000 565.440 ;
        RECT 3.990 555.920 596.000 564.040 ;
        RECT 3.990 554.520 595.600 555.920 ;
        RECT 3.990 547.760 596.000 554.520 ;
        RECT 4.400 546.360 596.000 547.760 ;
        RECT 3.990 538.240 596.000 546.360 ;
        RECT 3.990 536.840 595.600 538.240 ;
        RECT 3.990 530.080 596.000 536.840 ;
        RECT 4.400 528.680 596.000 530.080 ;
        RECT 3.990 520.560 596.000 528.680 ;
        RECT 3.990 519.160 595.600 520.560 ;
        RECT 3.990 512.400 596.000 519.160 ;
        RECT 4.400 511.000 596.000 512.400 ;
        RECT 3.990 502.880 596.000 511.000 ;
        RECT 3.990 501.480 595.600 502.880 ;
        RECT 3.990 494.720 596.000 501.480 ;
        RECT 4.400 493.320 596.000 494.720 ;
        RECT 3.990 485.200 596.000 493.320 ;
        RECT 3.990 483.800 595.600 485.200 ;
        RECT 3.990 477.040 596.000 483.800 ;
        RECT 4.400 475.640 596.000 477.040 ;
        RECT 3.990 467.520 596.000 475.640 ;
        RECT 3.990 466.120 595.600 467.520 ;
        RECT 3.990 459.360 596.000 466.120 ;
        RECT 4.400 457.960 596.000 459.360 ;
        RECT 3.990 449.840 596.000 457.960 ;
        RECT 3.990 448.440 595.600 449.840 ;
        RECT 3.990 441.680 596.000 448.440 ;
        RECT 4.400 440.280 596.000 441.680 ;
        RECT 3.990 432.160 596.000 440.280 ;
        RECT 3.990 430.760 595.600 432.160 ;
        RECT 3.990 424.000 596.000 430.760 ;
        RECT 4.400 422.600 596.000 424.000 ;
        RECT 3.990 414.480 596.000 422.600 ;
        RECT 3.990 413.080 595.600 414.480 ;
        RECT 3.990 406.320 596.000 413.080 ;
        RECT 4.400 404.920 596.000 406.320 ;
        RECT 3.990 396.800 596.000 404.920 ;
        RECT 3.990 395.400 595.600 396.800 ;
        RECT 3.990 388.640 596.000 395.400 ;
        RECT 4.400 387.240 596.000 388.640 ;
        RECT 3.990 379.120 596.000 387.240 ;
        RECT 3.990 377.720 595.600 379.120 ;
        RECT 3.990 370.960 596.000 377.720 ;
        RECT 4.400 369.560 596.000 370.960 ;
        RECT 3.990 361.440 596.000 369.560 ;
        RECT 3.990 360.040 595.600 361.440 ;
        RECT 3.990 353.280 596.000 360.040 ;
        RECT 4.400 351.880 596.000 353.280 ;
        RECT 3.990 343.760 596.000 351.880 ;
        RECT 3.990 342.360 595.600 343.760 ;
        RECT 3.990 335.600 596.000 342.360 ;
        RECT 4.400 334.200 596.000 335.600 ;
        RECT 3.990 326.080 596.000 334.200 ;
        RECT 3.990 324.680 595.600 326.080 ;
        RECT 3.990 317.920 596.000 324.680 ;
        RECT 4.400 316.520 596.000 317.920 ;
        RECT 3.990 308.400 596.000 316.520 ;
        RECT 3.990 307.000 595.600 308.400 ;
        RECT 3.990 300.240 596.000 307.000 ;
        RECT 4.400 298.840 596.000 300.240 ;
        RECT 3.990 290.720 596.000 298.840 ;
        RECT 3.990 289.320 595.600 290.720 ;
        RECT 3.990 282.560 596.000 289.320 ;
        RECT 4.400 281.160 596.000 282.560 ;
        RECT 3.990 273.040 596.000 281.160 ;
        RECT 3.990 271.640 595.600 273.040 ;
        RECT 3.990 264.880 596.000 271.640 ;
        RECT 4.400 263.480 596.000 264.880 ;
        RECT 3.990 255.360 596.000 263.480 ;
        RECT 3.990 253.960 595.600 255.360 ;
        RECT 3.990 247.200 596.000 253.960 ;
        RECT 4.400 245.800 596.000 247.200 ;
        RECT 3.990 237.680 596.000 245.800 ;
        RECT 3.990 236.280 595.600 237.680 ;
        RECT 3.990 229.520 596.000 236.280 ;
        RECT 4.400 228.120 596.000 229.520 ;
        RECT 3.990 220.000 596.000 228.120 ;
        RECT 3.990 218.600 595.600 220.000 ;
        RECT 3.990 211.840 596.000 218.600 ;
        RECT 4.400 210.440 596.000 211.840 ;
        RECT 3.990 202.320 596.000 210.440 ;
        RECT 3.990 200.920 595.600 202.320 ;
        RECT 3.990 194.160 596.000 200.920 ;
        RECT 4.400 192.760 596.000 194.160 ;
        RECT 3.990 184.640 596.000 192.760 ;
        RECT 3.990 183.240 595.600 184.640 ;
        RECT 3.990 176.480 596.000 183.240 ;
        RECT 4.400 175.080 596.000 176.480 ;
        RECT 3.990 166.960 596.000 175.080 ;
        RECT 3.990 165.560 595.600 166.960 ;
        RECT 3.990 158.800 596.000 165.560 ;
        RECT 4.400 157.400 596.000 158.800 ;
        RECT 3.990 149.280 596.000 157.400 ;
        RECT 3.990 147.880 595.600 149.280 ;
        RECT 3.990 141.120 596.000 147.880 ;
        RECT 4.400 139.720 596.000 141.120 ;
        RECT 3.990 131.600 596.000 139.720 ;
        RECT 3.990 130.200 595.600 131.600 ;
        RECT 3.990 123.440 596.000 130.200 ;
        RECT 4.400 122.040 596.000 123.440 ;
        RECT 3.990 113.920 596.000 122.040 ;
        RECT 3.990 112.520 595.600 113.920 ;
        RECT 3.990 105.760 596.000 112.520 ;
        RECT 4.400 104.360 596.000 105.760 ;
        RECT 3.990 96.240 596.000 104.360 ;
        RECT 3.990 94.840 595.600 96.240 ;
        RECT 3.990 88.080 596.000 94.840 ;
        RECT 4.400 86.680 596.000 88.080 ;
        RECT 3.990 78.560 596.000 86.680 ;
        RECT 3.990 77.160 595.600 78.560 ;
        RECT 3.990 70.400 596.000 77.160 ;
        RECT 4.400 69.000 596.000 70.400 ;
        RECT 3.990 60.880 596.000 69.000 ;
        RECT 3.990 59.480 595.600 60.880 ;
        RECT 3.990 52.720 596.000 59.480 ;
        RECT 4.400 51.320 596.000 52.720 ;
        RECT 3.990 43.200 596.000 51.320 ;
        RECT 3.990 41.800 595.600 43.200 ;
        RECT 3.990 35.040 596.000 41.800 ;
        RECT 4.400 33.640 596.000 35.040 ;
        RECT 3.990 25.520 596.000 33.640 ;
        RECT 3.990 24.120 595.600 25.520 ;
        RECT 3.990 17.360 596.000 24.120 ;
        RECT 4.400 15.960 596.000 17.360 ;
        RECT 3.990 10.715 596.000 15.960 ;
      LAYER met4 ;
        RECT 80.335 13.095 120.640 476.505 ;
        RECT 123.040 13.095 123.940 476.505 ;
        RECT 126.340 13.095 170.640 476.505 ;
        RECT 173.040 13.095 173.940 476.505 ;
        RECT 176.340 13.095 220.640 476.505 ;
        RECT 223.040 13.095 223.940 476.505 ;
        RECT 226.340 13.095 270.640 476.505 ;
        RECT 273.040 13.095 273.940 476.505 ;
        RECT 276.340 13.095 320.640 476.505 ;
        RECT 323.040 13.095 323.940 476.505 ;
        RECT 326.340 13.095 370.640 476.505 ;
        RECT 373.040 13.095 373.940 476.505 ;
        RECT 376.340 13.095 420.640 476.505 ;
        RECT 423.040 13.095 423.940 476.505 ;
        RECT 426.340 13.095 470.640 476.505 ;
        RECT 473.040 13.095 473.940 476.505 ;
        RECT 476.340 13.095 519.505 476.505 ;
      LAYER met5 ;
        RECT 236.100 266.100 283.700 267.700 ;
  END
END pipelined_mult
END LIBRARY

