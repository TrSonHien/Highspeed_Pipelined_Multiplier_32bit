VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pipelined_mult
  CLASS BLOCK ;
  FOREIGN pipelined_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.340 10.640 95.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.340 10.640 165.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.340 10.640 235.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.340 10.640 305.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.340 10.640 375.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 444.340 10.640 445.940 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.340 10.640 515.940 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 544.420 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 100.030 544.420 101.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 170.030 544.420 171.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 240.030 544.420 241.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 310.030 544.420 311.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 380.030 544.420 381.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 450.030 544.420 451.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 520.030 544.420 521.630 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.040 10.640 92.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.040 10.640 162.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 231.040 10.640 232.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.040 10.640 302.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 441.040 10.640 442.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 511.040 10.640 512.640 538.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 544.420 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 96.730 544.420 98.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 166.730 544.420 168.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 236.730 544.420 238.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 306.730 544.420 308.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 376.730 544.420 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 446.730 544.420 448.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 516.730 544.420 518.330 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END a[9]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END b[0]
  PIN b[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 291.270 0.000 291.550 4.000 ;
    END
  END b[10]
  PIN b[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END b[11]
  PIN b[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END b[12]
  PIN b[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END b[13]
  PIN b[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END b[14]
  PIN b[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 374.070 0.000 374.350 4.000 ;
    END
  END b[15]
  PIN b[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END b[16]
  PIN b[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END b[17]
  PIN b[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END b[18]
  PIN b[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END b[19]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END b[1]
  PIN b[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END b[20]
  PIN b[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END b[21]
  PIN b[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END b[22]
  PIN b[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END b[23]
  PIN b[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END b[24]
  PIN b[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END b[25]
  PIN b[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END b[26]
  PIN b[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END b[27]
  PIN b[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END b[28]
  PIN b[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END b[29]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END b[2]
  PIN b[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END b[30]
  PIN b[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END b[31]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END b[7]
  PIN b[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END b[8]
  PIN b[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END b[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END clk
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 380.840 550.000 381.440 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 217.640 550.000 218.240 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 233.960 550.000 234.560 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 250.280 550.000 250.880 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 266.600 550.000 267.200 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 282.920 550.000 283.520 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 299.240 550.000 299.840 ;
    END
  END p[15]
  PIN p[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 315.560 550.000 316.160 ;
    END
  END p[16]
  PIN p[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 331.880 550.000 332.480 ;
    END
  END p[17]
  PIN p[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 348.200 550.000 348.800 ;
    END
  END p[18]
  PIN p[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 364.520 550.000 365.120 ;
    END
  END p[19]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 397.160 550.000 397.760 ;
    END
  END p[1]
  PIN p[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 54.440 550.000 55.040 ;
    END
  END p[20]
  PIN p[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 70.760 550.000 71.360 ;
    END
  END p[21]
  PIN p[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 87.080 550.000 87.680 ;
    END
  END p[22]
  PIN p[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 103.400 550.000 104.000 ;
    END
  END p[23]
  PIN p[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 119.720 550.000 120.320 ;
    END
  END p[24]
  PIN p[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 136.040 550.000 136.640 ;
    END
  END p[25]
  PIN p[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 152.360 550.000 152.960 ;
    END
  END p[26]
  PIN p[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 168.680 550.000 169.280 ;
    END
  END p[27]
  PIN p[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 185.000 550.000 185.600 ;
    END
  END p[28]
  PIN p[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 201.320 550.000 201.920 ;
    END
  END p[29]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 413.480 550.000 414.080 ;
    END
  END p[2]
  PIN p[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 21.800 550.000 22.400 ;
    END
  END p[30]
  PIN p[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 38.120 550.000 38.720 ;
    END
  END p[31]
  PIN p[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 419.610 546.000 419.890 550.000 ;
    END
  END p[32]
  PIN p[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 436.630 546.000 436.910 550.000 ;
    END
  END p[33]
  PIN p[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 453.650 546.000 453.930 550.000 ;
    END
  END p[34]
  PIN p[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 470.670 546.000 470.950 550.000 ;
    END
  END p[35]
  PIN p[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 487.690 546.000 487.970 550.000 ;
    END
  END p[36]
  PIN p[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 504.710 546.000 504.990 550.000 ;
    END
  END p[37]
  PIN p[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 521.730 546.000 522.010 550.000 ;
    END
  END p[38]
  PIN p[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 538.750 546.000 539.030 550.000 ;
    END
  END p[39]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 429.800 550.000 430.400 ;
    END
  END p[3]
  PIN p[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 249.410 546.000 249.690 550.000 ;
    END
  END p[40]
  PIN p[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 266.430 546.000 266.710 550.000 ;
    END
  END p[41]
  PIN p[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 283.450 546.000 283.730 550.000 ;
    END
  END p[42]
  PIN p[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 300.470 546.000 300.750 550.000 ;
    END
  END p[43]
  PIN p[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.490 546.000 317.770 550.000 ;
    END
  END p[44]
  PIN p[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 334.510 546.000 334.790 550.000 ;
    END
  END p[45]
  PIN p[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 351.530 546.000 351.810 550.000 ;
    END
  END p[46]
  PIN p[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 368.550 546.000 368.830 550.000 ;
    END
  END p[47]
  PIN p[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 385.570 546.000 385.850 550.000 ;
    END
  END p[48]
  PIN p[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 402.590 546.000 402.870 550.000 ;
    END
  END p[49]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 446.120 550.000 446.720 ;
    END
  END p[4]
  PIN p[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.210 546.000 79.490 550.000 ;
    END
  END p[50]
  PIN p[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 546.000 96.510 550.000 ;
    END
  END p[51]
  PIN p[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.250 546.000 113.530 550.000 ;
    END
  END p[52]
  PIN p[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.270 546.000 130.550 550.000 ;
    END
  END p[53]
  PIN p[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 147.290 546.000 147.570 550.000 ;
    END
  END p[54]
  PIN p[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 546.000 164.590 550.000 ;
    END
  END p[55]
  PIN p[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 181.330 546.000 181.610 550.000 ;
    END
  END p[56]
  PIN p[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 546.000 198.630 550.000 ;
    END
  END p[57]
  PIN p[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.370 546.000 215.650 550.000 ;
    END
  END p[58]
  PIN p[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 232.390 546.000 232.670 550.000 ;
    END
  END p[59]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 462.440 550.000 463.040 ;
    END
  END p[5]
  PIN p[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 11.130 546.000 11.410 550.000 ;
    END
  END p[60]
  PIN p[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.150 546.000 28.430 550.000 ;
    END
  END p[61]
  PIN p[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 546.000 45.450 550.000 ;
    END
  END p[62]
  PIN p[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 62.190 546.000 62.470 550.000 ;
    END
  END p[63]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 478.760 550.000 479.360 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 495.080 550.000 495.680 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 511.400 550.000 512.000 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 527.720 550.000 528.320 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 544.370 538.645 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 4.210 10.640 544.480 538.800 ;
      LAYER met2 ;
        RECT 4.230 545.720 10.850 546.000 ;
        RECT 11.690 545.720 27.870 546.000 ;
        RECT 28.710 545.720 44.890 546.000 ;
        RECT 45.730 545.720 61.910 546.000 ;
        RECT 62.750 545.720 78.930 546.000 ;
        RECT 79.770 545.720 95.950 546.000 ;
        RECT 96.790 545.720 112.970 546.000 ;
        RECT 113.810 545.720 129.990 546.000 ;
        RECT 130.830 545.720 147.010 546.000 ;
        RECT 147.850 545.720 164.030 546.000 ;
        RECT 164.870 545.720 181.050 546.000 ;
        RECT 181.890 545.720 198.070 546.000 ;
        RECT 198.910 545.720 215.090 546.000 ;
        RECT 215.930 545.720 232.110 546.000 ;
        RECT 232.950 545.720 249.130 546.000 ;
        RECT 249.970 545.720 266.150 546.000 ;
        RECT 266.990 545.720 283.170 546.000 ;
        RECT 284.010 545.720 300.190 546.000 ;
        RECT 301.030 545.720 317.210 546.000 ;
        RECT 318.050 545.720 334.230 546.000 ;
        RECT 335.070 545.720 351.250 546.000 ;
        RECT 352.090 545.720 368.270 546.000 ;
        RECT 369.110 545.720 385.290 546.000 ;
        RECT 386.130 545.720 402.310 546.000 ;
        RECT 403.150 545.720 419.330 546.000 ;
        RECT 420.170 545.720 436.350 546.000 ;
        RECT 437.190 545.720 453.370 546.000 ;
        RECT 454.210 545.720 470.390 546.000 ;
        RECT 471.230 545.720 487.410 546.000 ;
        RECT 488.250 545.720 504.430 546.000 ;
        RECT 505.270 545.720 521.450 546.000 ;
        RECT 522.290 545.720 538.470 546.000 ;
        RECT 539.310 545.720 543.620 546.000 ;
        RECT 4.230 4.280 543.620 545.720 ;
        RECT 4.230 4.000 9.470 4.280 ;
        RECT 10.310 4.000 26.030 4.280 ;
        RECT 26.870 4.000 42.590 4.280 ;
        RECT 43.430 4.000 59.150 4.280 ;
        RECT 59.990 4.000 75.710 4.280 ;
        RECT 76.550 4.000 92.270 4.280 ;
        RECT 93.110 4.000 108.830 4.280 ;
        RECT 109.670 4.000 125.390 4.280 ;
        RECT 126.230 4.000 141.950 4.280 ;
        RECT 142.790 4.000 158.510 4.280 ;
        RECT 159.350 4.000 175.070 4.280 ;
        RECT 175.910 4.000 191.630 4.280 ;
        RECT 192.470 4.000 208.190 4.280 ;
        RECT 209.030 4.000 224.750 4.280 ;
        RECT 225.590 4.000 241.310 4.280 ;
        RECT 242.150 4.000 257.870 4.280 ;
        RECT 258.710 4.000 274.430 4.280 ;
        RECT 275.270 4.000 290.990 4.280 ;
        RECT 291.830 4.000 307.550 4.280 ;
        RECT 308.390 4.000 324.110 4.280 ;
        RECT 324.950 4.000 340.670 4.280 ;
        RECT 341.510 4.000 357.230 4.280 ;
        RECT 358.070 4.000 373.790 4.280 ;
        RECT 374.630 4.000 390.350 4.280 ;
        RECT 391.190 4.000 406.910 4.280 ;
        RECT 407.750 4.000 423.470 4.280 ;
        RECT 424.310 4.000 440.030 4.280 ;
        RECT 440.870 4.000 456.590 4.280 ;
        RECT 457.430 4.000 473.150 4.280 ;
        RECT 473.990 4.000 489.710 4.280 ;
        RECT 490.550 4.000 506.270 4.280 ;
        RECT 507.110 4.000 522.830 4.280 ;
        RECT 523.670 4.000 539.390 4.280 ;
        RECT 540.230 4.000 543.620 4.280 ;
      LAYER met3 ;
        RECT 3.990 536.880 546.000 538.725 ;
        RECT 4.400 535.480 546.000 536.880 ;
        RECT 3.990 528.720 546.000 535.480 ;
        RECT 3.990 527.320 545.600 528.720 ;
        RECT 3.990 520.560 546.000 527.320 ;
        RECT 4.400 519.160 546.000 520.560 ;
        RECT 3.990 512.400 546.000 519.160 ;
        RECT 3.990 511.000 545.600 512.400 ;
        RECT 3.990 504.240 546.000 511.000 ;
        RECT 4.400 502.840 546.000 504.240 ;
        RECT 3.990 496.080 546.000 502.840 ;
        RECT 3.990 494.680 545.600 496.080 ;
        RECT 3.990 487.920 546.000 494.680 ;
        RECT 4.400 486.520 546.000 487.920 ;
        RECT 3.990 479.760 546.000 486.520 ;
        RECT 3.990 478.360 545.600 479.760 ;
        RECT 3.990 471.600 546.000 478.360 ;
        RECT 4.400 470.200 546.000 471.600 ;
        RECT 3.990 463.440 546.000 470.200 ;
        RECT 3.990 462.040 545.600 463.440 ;
        RECT 3.990 455.280 546.000 462.040 ;
        RECT 4.400 453.880 546.000 455.280 ;
        RECT 3.990 447.120 546.000 453.880 ;
        RECT 3.990 445.720 545.600 447.120 ;
        RECT 3.990 438.960 546.000 445.720 ;
        RECT 4.400 437.560 546.000 438.960 ;
        RECT 3.990 430.800 546.000 437.560 ;
        RECT 3.990 429.400 545.600 430.800 ;
        RECT 3.990 422.640 546.000 429.400 ;
        RECT 4.400 421.240 546.000 422.640 ;
        RECT 3.990 414.480 546.000 421.240 ;
        RECT 3.990 413.080 545.600 414.480 ;
        RECT 3.990 406.320 546.000 413.080 ;
        RECT 4.400 404.920 546.000 406.320 ;
        RECT 3.990 398.160 546.000 404.920 ;
        RECT 3.990 396.760 545.600 398.160 ;
        RECT 3.990 390.000 546.000 396.760 ;
        RECT 4.400 388.600 546.000 390.000 ;
        RECT 3.990 381.840 546.000 388.600 ;
        RECT 3.990 380.440 545.600 381.840 ;
        RECT 3.990 373.680 546.000 380.440 ;
        RECT 4.400 372.280 546.000 373.680 ;
        RECT 3.990 365.520 546.000 372.280 ;
        RECT 3.990 364.120 545.600 365.520 ;
        RECT 3.990 357.360 546.000 364.120 ;
        RECT 4.400 355.960 546.000 357.360 ;
        RECT 3.990 349.200 546.000 355.960 ;
        RECT 3.990 347.800 545.600 349.200 ;
        RECT 3.990 341.040 546.000 347.800 ;
        RECT 4.400 339.640 546.000 341.040 ;
        RECT 3.990 332.880 546.000 339.640 ;
        RECT 3.990 331.480 545.600 332.880 ;
        RECT 3.990 324.720 546.000 331.480 ;
        RECT 4.400 323.320 546.000 324.720 ;
        RECT 3.990 316.560 546.000 323.320 ;
        RECT 3.990 315.160 545.600 316.560 ;
        RECT 3.990 308.400 546.000 315.160 ;
        RECT 4.400 307.000 546.000 308.400 ;
        RECT 3.990 300.240 546.000 307.000 ;
        RECT 3.990 298.840 545.600 300.240 ;
        RECT 3.990 292.080 546.000 298.840 ;
        RECT 4.400 290.680 546.000 292.080 ;
        RECT 3.990 283.920 546.000 290.680 ;
        RECT 3.990 282.520 545.600 283.920 ;
        RECT 3.990 275.760 546.000 282.520 ;
        RECT 4.400 274.360 546.000 275.760 ;
        RECT 3.990 267.600 546.000 274.360 ;
        RECT 3.990 266.200 545.600 267.600 ;
        RECT 3.990 259.440 546.000 266.200 ;
        RECT 4.400 258.040 546.000 259.440 ;
        RECT 3.990 251.280 546.000 258.040 ;
        RECT 3.990 249.880 545.600 251.280 ;
        RECT 3.990 243.120 546.000 249.880 ;
        RECT 4.400 241.720 546.000 243.120 ;
        RECT 3.990 234.960 546.000 241.720 ;
        RECT 3.990 233.560 545.600 234.960 ;
        RECT 3.990 226.800 546.000 233.560 ;
        RECT 4.400 225.400 546.000 226.800 ;
        RECT 3.990 218.640 546.000 225.400 ;
        RECT 3.990 217.240 545.600 218.640 ;
        RECT 3.990 210.480 546.000 217.240 ;
        RECT 4.400 209.080 546.000 210.480 ;
        RECT 3.990 202.320 546.000 209.080 ;
        RECT 3.990 200.920 545.600 202.320 ;
        RECT 3.990 194.160 546.000 200.920 ;
        RECT 4.400 192.760 546.000 194.160 ;
        RECT 3.990 186.000 546.000 192.760 ;
        RECT 3.990 184.600 545.600 186.000 ;
        RECT 3.990 177.840 546.000 184.600 ;
        RECT 4.400 176.440 546.000 177.840 ;
        RECT 3.990 169.680 546.000 176.440 ;
        RECT 3.990 168.280 545.600 169.680 ;
        RECT 3.990 161.520 546.000 168.280 ;
        RECT 4.400 160.120 546.000 161.520 ;
        RECT 3.990 153.360 546.000 160.120 ;
        RECT 3.990 151.960 545.600 153.360 ;
        RECT 3.990 145.200 546.000 151.960 ;
        RECT 4.400 143.800 546.000 145.200 ;
        RECT 3.990 137.040 546.000 143.800 ;
        RECT 3.990 135.640 545.600 137.040 ;
        RECT 3.990 128.880 546.000 135.640 ;
        RECT 4.400 127.480 546.000 128.880 ;
        RECT 3.990 120.720 546.000 127.480 ;
        RECT 3.990 119.320 545.600 120.720 ;
        RECT 3.990 112.560 546.000 119.320 ;
        RECT 4.400 111.160 546.000 112.560 ;
        RECT 3.990 104.400 546.000 111.160 ;
        RECT 3.990 103.000 545.600 104.400 ;
        RECT 3.990 96.240 546.000 103.000 ;
        RECT 4.400 94.840 546.000 96.240 ;
        RECT 3.990 88.080 546.000 94.840 ;
        RECT 3.990 86.680 545.600 88.080 ;
        RECT 3.990 79.920 546.000 86.680 ;
        RECT 4.400 78.520 546.000 79.920 ;
        RECT 3.990 71.760 546.000 78.520 ;
        RECT 3.990 70.360 545.600 71.760 ;
        RECT 3.990 63.600 546.000 70.360 ;
        RECT 4.400 62.200 546.000 63.600 ;
        RECT 3.990 55.440 546.000 62.200 ;
        RECT 3.990 54.040 545.600 55.440 ;
        RECT 3.990 47.280 546.000 54.040 ;
        RECT 4.400 45.880 546.000 47.280 ;
        RECT 3.990 39.120 546.000 45.880 ;
        RECT 3.990 37.720 545.600 39.120 ;
        RECT 3.990 30.960 546.000 37.720 ;
        RECT 4.400 29.560 546.000 30.960 ;
        RECT 3.990 22.800 546.000 29.560 ;
        RECT 3.990 21.400 545.600 22.800 ;
        RECT 3.990 14.640 546.000 21.400 ;
        RECT 4.400 13.240 546.000 14.640 ;
        RECT 3.990 10.715 546.000 13.240 ;
      LAYER met4 ;
        RECT 49.975 13.095 90.640 476.505 ;
        RECT 93.040 13.095 93.940 476.505 ;
        RECT 96.340 13.095 160.640 476.505 ;
        RECT 163.040 13.095 163.940 476.505 ;
        RECT 166.340 13.095 230.640 476.505 ;
        RECT 233.040 13.095 233.940 476.505 ;
        RECT 236.340 13.095 300.640 476.505 ;
        RECT 303.040 13.095 303.940 476.505 ;
        RECT 306.340 13.095 370.640 476.505 ;
        RECT 373.040 13.095 373.940 476.505 ;
        RECT 376.340 13.095 440.640 476.505 ;
        RECT 443.040 13.095 443.940 476.505 ;
        RECT 446.340 13.095 505.705 476.505 ;
  END
END pipelined_mult
END LIBRARY

