* NGSPICE file created from pipelined_mult.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

.subckt pipelined_mult VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16] a[17]
+ a[18] a[19] a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29] a[2]
+ a[30] a[31] a[3] a[4] a[5] a[6] a[7] a[8] a[9] b[0] b[10] b[11] b[12] b[13] b[14]
+ b[15] b[16] b[17] b[18] b[19] b[1] b[20] b[21] b[22] b[23] b[24] b[25] b[26] b[27]
+ b[28] b[29] b[2] b[30] b[31] b[3] b[4] b[5] b[6] b[7] b[8] b[9] clk p[0] p[10] p[11]
+ p[12] p[13] p[14] p[15] p[16] p[17] p[18] p[19] p[1] p[20] p[21] p[22] p[23] p[24]
+ p[25] p[26] p[27] p[28] p[29] p[2] p[30] p[31] p[32] p[33] p[34] p[35] p[36] p[37]
+ p[38] p[39] p[3] p[40] p[41] p[42] p[43] p[44] p[45] p[46] p[47] p[48] p[49] p[4]
+ p[50] p[51] p[52] p[53] p[54] p[55] p[56] p[57] p[58] p[59] p[5] p[60] p[61] p[62]
+ p[63] p[6] p[7] p[8] p[9] rst
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit293 a_l\[4\] VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__buf_2
X_18869_ net413 _09748_ _09756_ _09758_ VGND VGND VPWR VPWR _09761_ sky130_fd_sc_hd__o211ai_4
Xsplit282 b_l\[9\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_38_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20762_ clknet_leaf_3_clk _00402_ VGND VGND VPWR VPWR a_h\[0\] sky130_fd_sc_hd__dfxtp_4
XFILLER_62_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20693_ clknet_leaf_4_clk _00333_ VGND VGND VPWR VPWR p_hl\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold362 p_ll\[19\] VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 p_hh_pipe\[4\] VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 term_low\[5\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold395 p_ll\[21\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20127_ _01218_ _01361_ _01362_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__o21a_1
XFILLER_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20058_ _01285_ _01286_ _09286_ _09362_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__o2bb2a_1
X_11900_ net682 net492 VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__nand2_2
X_12880_ net396 _03756_ _03755_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a21o_1
X_11831_ _02766_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__nor2_1
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14550_ _05451_ _05439_ _05450_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__nand3_4
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11762_ net979 _02641_ _02643_ _02644_ _02664_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__a32oi_2
X_13501_ _02082_ _04134_ _04350_ _04348_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__o22a_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11693_ _09460_ _09602_ net462 _02629_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__o22a_1
X_10713_ p_hl\[14\] p_lh\[14\] VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__xor2_1
X_14481_ _05383_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__inv_2
X_16220_ net570 net541 VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__nand2_1
X_10644_ _01686_ _01687_ _01680_ _01684_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__o211a_1
X_13432_ _09220_ _09406_ _04338_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_24_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16151_ net841 net496 net491 net629 VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__a22oi_2
X_13363_ net763 net705 _04272_ _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__a22oi_2
XFILLER_10_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10575_ _09690_ net1339 VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__and2_1
X_12314_ _03242_ _03245_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__nand2_1
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer7 net800 VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_58_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15102_ net751 net745 net640 net635 VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__and4_4
X_16082_ net607 net512 VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__nand2_1
X_13294_ _04205_ _04157_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__nand2_1
XFILLER_6_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12245_ _03043_ net483 net687 a_h\[3\] net475 VGND VGND VPWR VPWR _03179_ sky130_fd_sc_hd__a32oi_2
XPHY_EDGE_ROW_2_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19910_ _01126_ _01129_ net589 net721 VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__and4_4
X_15033_ _05928_ _05930_ _09308_ _09482_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_39_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12176_ _03104_ _03106_ _03109_ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__nand3_1
XFILLER_123_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19841_ _01054_ _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__nand2_1
X_11127_ net691 net967 net525 net1052 _02063_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__a41o_1
X_16984_ _07620_ _07622_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__nand2_1
XFILLER_110_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19772_ net877 net548 VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__nand2_1
X_15935_ _06806_ _06811_ _06810_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__a21oi_1
X_11058_ _01959_ _01963_ _01961_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__a21boi_1
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18723_ net619 net887 net1082 net737 VGND VGND VPWR VPWR _09608_ sky130_fd_sc_hd__nand4_1
X_15866_ _06655_ _06662_ _06663_ _06667_ _06578_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__a32oi_4
XFILLER_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18654_ net626 net732 VGND VGND VPWR VPWR _09533_ sky130_fd_sc_hd__nand2_2
XFILLER_37_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17605_ _08413_ _08418_ VGND VGND VPWR VPWR _08469_ sky130_fd_sc_hd__nand2_1
X_18585_ _09199_ _09264_ net457 _06681_ _09454_ VGND VGND VPWR VPWR _09457_ sky130_fd_sc_hd__o221ai_2
X_14817_ net736 net668 net663 net739 VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__a22oi_4
X_15797_ _06600_ _06607_ _06603_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__a21oi_1
X_17536_ _09297_ _09646_ _08396_ _08398_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__o22ai_2
XPHY_EDGE_ROW_48_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14748_ _05647_ _05642_ _05539_ _05507_ _05648_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__o2111ai_2
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17467_ _08328_ _08330_ _08301_ VGND VGND VPWR VPWR _08333_ sky130_fd_sc_hd__o21ai_1
X_14679_ net425 _05577_ net426 VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__a21oi_2
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16418_ _07187_ _07290_ _07291_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__nand3_2
X_17398_ _08261_ _08164_ _08260_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_43_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19206_ _10099_ _10084_ VGND VGND VPWR VPWR _10103_ sky130_fd_sc_hd__nand2_2
X_16349_ _07123_ _07126_ net280 _07149_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__a2bb2oi_1
X_19137_ _10026_ _10027_ VGND VGND VPWR VPWR _10028_ sky130_fd_sc_hd__nand2_1
X_19068_ _09925_ _09950_ _09952_ VGND VGND VPWR VPWR _09959_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_113_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18019_ net779 net615 VGND VGND VPWR VPWR _08869_ sky130_fd_sc_hd__nand2_1
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20745_ clknet_leaf_42_clk _00385_ VGND VGND VPWR VPWR p_ll\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20676_ clknet_leaf_55_clk _00316_ VGND VGND VPWR VPWR p_hl\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire517 net518 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_21_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10360_ net471 _01322_ net794 VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10291_ _00558_ _00579_ net797 VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__a21oi_1
X_12030_ _02965_ _02964_ net796 VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13981_ _04876_ _04883_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__o21ai_1
X_15720_ net966 net541 VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__nand2_1
XFILLER_74_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12932_ _03802_ _03803_ _03857_ net175 VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a22o_1
X_15651_ _06531_ _06515_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__nand2_1
XFILLER_74_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12863_ _03602_ _03705_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__or2_1
X_14602_ _05463_ _05464_ _05497_ _05498_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__nand4_1
XFILLER_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ net628 net522 VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__nand2_1
X_11814_ _02745_ _02746_ _02730_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__nand3_1
X_12794_ _03720_ _03716_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__nand2_1
X_18370_ _09124_ _09128_ _09219_ VGND VGND VPWR VPWR _09223_ sky130_fd_sc_hd__a21oi_4
X_11745_ _02677_ _02681_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__nand2_2
X_17321_ net341 _08184_ _08186_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__nand3_1
X_14533_ _05428_ _05430_ _05432_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__a21boi_1
X_17252_ _08100_ net450 _08098_ net342 _08116_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__o2111ai_4
X_14464_ _05362_ _05363_ _05219_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__a21o_1
X_16203_ net973 net484 VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__nand2_1
X_11676_ net646 net644 net546 net537 VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__nand4_1
X_13415_ net435 _04324_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_40_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10627_ p_hl\[0\] net1326 _01674_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__o21a_1
X_17183_ net571 net503 VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__nand2_1
X_14395_ _05168_ _05174_ _05294_ _05295_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__nand4_4
X_10558_ net793 net1267 VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__and2_1
XFILLER_127_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16134_ _06990_ _06994_ _07005_ _07007_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__o2bb2ai_1
X_13346_ _04215_ _04245_ _04247_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__o21a_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16065_ _06742_ _06827_ _06828_ _06728_ _06835_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__a32oi_1
XFILLER_108_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13277_ _04161_ _04165_ _04164_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__o21ai_1
XFILLER_52_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10489_ _01645_ term_high\[50\] term_high\[49\] net796 VGND VGND VPWR VPWR _01648_
+ sky130_fd_sc_hd__a31o_1
X_12228_ _03004_ _03022_ _03160_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__o21ai_4
X_15016_ _05911_ _05912_ VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__nor2_1
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12159_ _02852_ _03091_ _03092_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__nand3_1
XFILLER_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19824_ _00907_ _00908_ _00927_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__o21a_1
X_16967_ _07802_ _07804_ _07807_ _07829_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_68_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19755_ _00725_ _00727_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__and2_1
X_15918_ net617 net512 net505 net624 VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__a22o_1
XFILLER_83_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18706_ _09315_ _09320_ _09589_ VGND VGND VPWR VPWR _09590_ sky130_fd_sc_hd__o21ai_4
X_16898_ _07743_ _07745_ _07760_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__and3_1
XFILLER_92_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_56_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19686_ _00883_ _00885_ _00886_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__nand3_2
X_15849_ net191 _06652_ _06724_ _06725_ VGND VGND VPWR VPWR _06728_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_92_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18637_ _09513_ VGND VGND VPWR VPWR _09514_ sky130_fd_sc_hd__inv_2
XFILLER_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18568_ _09436_ _09437_ _09313_ VGND VGND VPWR VPWR _09440_ sky130_fd_sc_hd__a21oi_1
X_17519_ net941 net476 VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__and2_1
X_18499_ _09363_ _09357_ _09361_ VGND VGND VPWR VPWR _09364_ sky130_fd_sc_hd__a21o_1
XFILLER_33_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20530_ clknet_leaf_47_clk _00170_ VGND VGND VPWR VPWR term_low\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20461_ clknet_leaf_14_clk _00101_ VGND VGND VPWR VPWR term_high\[53\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20392_ clknet_leaf_37_clk net1317 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfxtp_1
XFILLER_114_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_108_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11530_ _02464_ _02466_ _02465_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__and3_1
XFILLER_24_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_83_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20728_ clknet_leaf_6_clk _00368_ VGND VGND VPWR VPWR p_lh\[30\] sky130_fd_sc_hd__dfxtp_1
Xwire303 _09346_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11461_ _02396_ _02399_ _02394_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__a21o_1
Xwire325 _02623_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__buf_6
X_20659_ clknet_leaf_10_clk _00299_ VGND VGND VPWR VPWR p_hh\[25\] sky130_fd_sc_hd__dfxtp_1
Xwire336 _09036_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10412_ _01574_ _01581_ _01582_ _01580_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__o31a_1
X_11392_ _02136_ net180 _02144_ _02234_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__o22ai_2
XFILLER_137_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13200_ _04120_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__inv_2
X_14180_ _05082_ net210 _04967_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13131_ _04053_ _04054_ _09504_ _09679_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__a211o_1
X_10343_ _01139_ VGND VGND VPWR VPWR _01150_ sky130_fd_sc_hd__inv_2
X_13062_ _03931_ _03932_ _03986_ _03987_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__a22o_1
X_10274_ term_low\[18\] term_mid\[18\] VGND VGND VPWR VPWR _10137_ sky130_fd_sc_hd__and2_1
XFILLER_3_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12013_ _02936_ _02937_ _02946_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_92_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17870_ _08726_ _08727_ _09319_ _09679_ VGND VGND VPWR VPWR _08730_ sky130_fd_sc_hd__o2bb2a_1
X_16821_ _07664_ net278 _07688_ _07689_ VGND VGND VPWR VPWR _07692_ sky130_fd_sc_hd__o2bb2ai_1
X_16752_ _07478_ _07467_ _07469_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__o21ai_1
XFILLER_120_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone226 b_h\[4\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__clkbuf_16
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19540_ _09220_ _09373_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__nor2_1
X_15703_ _06578_ _06579_ _06580_ _06538_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__o22a_2
XFILLER_65_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13964_ net318 _04761_ _04763_ _04727_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__a31oi_2
X_16683_ _07491_ _07549_ _07551_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__nand3_2
X_12915_ _03839_ _03840_ _03732_ VGND VGND VPWR VPWR _03843_ sky130_fd_sc_hd__a21oi_1
XFILLER_46_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13895_ _04797_ _04798_ _04667_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19471_ _09264_ _09286_ _00455_ _00653_ _00652_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__o221ai_4
X_15634_ _06475_ _06478_ _06481_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__o21ai_2
X_12846_ _03772_ _03773_ _03727_ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_66_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18422_ net457 _06521_ net1100 net1148 _09274_ VGND VGND VPWR VPWR _09280_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_66_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _06444_ _06446_ net423 VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__a21oi_1
X_18353_ net1042 VGND VGND VPWR VPWR _09205_ sky130_fd_sc_hd__inv_2
XFILLER_15_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12777_ _03600_ _03609_ _03705_ net65 VGND VGND VPWR VPWR _03707_ sky130_fd_sc_hd__a31o_1
X_17304_ net573 net569 net498 net493 VGND VGND VPWR VPWR _08171_ sky130_fd_sc_hd__nand4_2
XFILLER_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14516_ net746 net668 VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__nand2_1
X_11728_ _02644_ _02664_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__nand2_1
X_18284_ _09028_ _09030_ _09124_ _09125_ VGND VGND VPWR VPWR _09130_ sky130_fd_sc_hd__a22o_1
X_15496_ _06364_ _06366_ _06384_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__o21bai_1
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11659_ _02585_ _02586_ _02592_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__nand3_2
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17235_ _07954_ _07951_ _07955_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__a21boi_1
X_14447_ _05346_ _05348_ _09308_ _09428_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__o2bb2ai_1
X_17166_ _07978_ _07984_ VGND VGND VPWR VPWR _08034_ sky130_fd_sc_hd__nand2_1
Xmax_cap603 net604 VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__buf_12
X_14378_ _02613_ net805 net761 net655 _05274_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__o2111ai_4
Xmax_cap625 a_l\[2\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__buf_8
X_16117_ _06992_ _06978_ _06991_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__and3_1
X_13329_ _04233_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nand2_1
Xmax_cap636 a_h\[15\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__buf_8
XFILLER_115_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap658 net661 VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__buf_12
X_17097_ net612 net476 VGND VGND VPWR VPWR _07966_ sky130_fd_sc_hd__nand2_1
Xmax_cap647 net648 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap669 a_h\[9\] VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__buf_12
X_16048_ _06787_ _06817_ _06922_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__a22oi_4
XFILLER_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19807_ b_l\[10\] net563 VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__nand2_2
XFILLER_29_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17999_ _08825_ net774 net632 VGND VGND VPWR VPWR _08850_ sky130_fd_sc_hd__nand3_1
X_19738_ _00810_ _00941_ _00939_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__o21ai_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19669_ net819 net552 VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__nand2_2
XFILLER_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20513_ clknet_leaf_31_clk _00153_ VGND VGND VPWR VPWR term_low\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20444_ clknet_leaf_27_clk _00084_ VGND VGND VPWR VPWR term_high\[36\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20375_ clknet_leaf_52_clk _00015_ VGND VGND VPWR VPWR b_l\[15\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_128_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10961_ net712 net517 VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__nand2_1
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12700_ _03629_ net475 net680 _03628_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__and4_1
X_13680_ _04516_ _04534_ _04530_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__a21boi_4
XFILLER_44_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12631_ _03559_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10892_ net794 net1205 VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__and2_1
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12562_ _03488_ _03489_ _03490_ VGND VGND VPWR VPWR _03494_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_61_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _06179_ _06186_ _06242_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__a21o_1
XFILLER_12_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11513_ net708 net487 VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__nand2_1
X_12493_ net1049 b_h\[4\] _03419_ _03423_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_61_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _06157_ _06175_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__nand2_1
X_14301_ net736 net690 net685 net740 VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a22oi_1
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire133 _00353_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
X_17020_ _07766_ _07772_ VGND VGND VPWR VPWR _07889_ sky130_fd_sc_hd__nand2_1
X_11444_ _02378_ _02380_ _02367_ _02371_ _02370_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__o221ai_4
Xwire155 _06298_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__buf_1
X_14232_ _05121_ _05131_ _05133_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__nand3_2
XFILLER_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11375_ _02312_ _02251_ _02311_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__nand3_4
X_14163_ _05067_ _05050_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__nand2_1
XFILLER_124_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13114_ _04036_ _04037_ _04033_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a21oi_1
X_18971_ _09730_ _09735_ _09862_ VGND VGND VPWR VPWR _09863_ sky130_fd_sc_hd__a21oi_1
X_10326_ term_low\[26\] term_mid\[26\] VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__nor2_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14094_ _04990_ _04993_ _04997_ net392 VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__o211ai_2
XFILLER_140_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17922_ net555 net473 VGND VGND VPWR VPWR _08780_ sky130_fd_sc_hd__nand2_1
X_10257_ net794 net1206 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__and2_1
X_13045_ _03969_ _03968_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__nand2_1
XFILLER_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17853_ _08613_ _08668_ _08667_ VGND VGND VPWR VPWR _08714_ sky130_fd_sc_hd__a21oi_1
X_10188_ net597 VGND VGND VPWR VPWR _09231_ sky130_fd_sc_hd__inv_12
XFILLER_38_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16804_ _07495_ _07671_ net590 net503 _07670_ VGND VGND VPWR VPWR _07675_ sky130_fd_sc_hd__o2111ai_2
X_17784_ _08643_ _08644_ VGND VGND VPWR VPWR _08646_ sky130_fd_sc_hd__xnor2_1
X_14996_ _05792_ _05865_ _05871_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__o21ai_1
X_16735_ net600 net594 net498 net493 VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__nand4_1
X_19523_ _00707_ _00708_ _00714_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13947_ _04779_ _04782_ _04843_ _04852_ _04784_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__o221ai_4
X_16666_ _07533_ _07535_ _07521_ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__nand3_4
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19454_ _00636_ _00639_ _00638_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__and3_1
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15617_ _06497_ _06498_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__nand2_2
X_18405_ _09243_ _09247_ _09257_ _09258_ VGND VGND VPWR VPWR _09261_ sky130_fd_sc_hd__o2bb2ai_1
X_13878_ _04783_ _04784_ net731 net709 VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__nand4_1
X_16597_ _07461_ _07462_ _07465_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__nand3_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12829_ _03739_ _03740_ _03756_ VGND VGND VPWR VPWR _03758_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19385_ _00561_ _00562_ _00563_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__nand3_1
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15548_ net611 net1041 VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__nand2_1
X_18336_ _09182_ _09185_ VGND VGND VPWR VPWR _09186_ sky130_fd_sc_hd__nand2_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18267_ net457 _06441_ _09030_ VGND VGND VPWR VPWR _09113_ sky130_fd_sc_hd__o21ai_2
XFILLER_30_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15479_ net719 net635 VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_96_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17218_ _08079_ _08082_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__nand2_1
X_18198_ _09040_ _09043_ VGND VGND VPWR VPWR _09045_ sky130_fd_sc_hd__nand2_1
Xmax_cap411 _09745_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_2
Xmax_cap422 _07030_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_2
X_17149_ _08009_ _08011_ _08013_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__nand3_1
Xmax_cap433 _04418_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__buf_1
Xmax_cap444 _01450_ VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap466 _01908_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_4
XFILLER_104_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap477 net478 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_8
Xmax_cap455 _05044_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_12
X_20160_ _01395_ _01396_ _01357_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__a21o_1
XFILLER_131_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap488 net490 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_6
Xmax_cap499 net500 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_12
X_20091_ _01209_ _01212_ net270 _01247_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__o22ai_4
XFILLER_84_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20427_ clknet_leaf_15_clk _00067_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfxtp_1
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11160_ _02019_ _02023_ _02021_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__a21oi_2
X_20358_ net794 net56 VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__and2_1
X_11091_ _02029_ _01999_ _02030_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__nand3_4
X_20289_ _01505_ _01506_ _01535_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14850_ _05746_ _05747_ _05669_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__a21oi_2
X_14781_ net756 net642 VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__nand2_2
X_13801_ net757 net683 VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__nand2_4
X_11993_ _02925_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__nand2_1
X_16520_ net572 net876 net544 net523 VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__and4_1
XFILLER_56_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13732_ _09264_ _09406_ _04490_ _04635_ _04634_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__o221ai_4
X_10944_ _01886_ _01887_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__nand2_1
XFILLER_44_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16451_ _07322_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__nand2_2
X_10875_ _09690_ net1239 VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__and2_1
X_13663_ _04552_ _04567_ _04566_ _04569_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__o211a_4
XFILLER_43_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16382_ _07225_ _07254_ _07255_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__nand3_2
X_12614_ _03539_ _03541_ _03536_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__a21o_1
X_13594_ _04500_ _04501_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__o21ai_4
X_15402_ _06246_ net1019 net715 _06243_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__a31o_1
XFILLER_43_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19170_ _10030_ _10031_ _10059_ VGND VGND VPWR VPWR _10064_ sky130_fd_sc_hd__nand3_2
X_12545_ _03473_ _03475_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__nand2_1
X_18121_ _08967_ _08966_ VGND VGND VPWR VPWR _08969_ sky130_fd_sc_hd__nand2_4
X_15333_ _06161_ _06165_ _06163_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__o21ai_1
XFILLER_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18052_ _08876_ _08867_ _08875_ _08864_ _08863_ VGND VGND VPWR VPWR _08901_ sky130_fd_sc_hd__a32oi_1
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17003_ _07708_ _07706_ _07707_ _07868_ _07869_ VGND VGND VPWR VPWR _07873_ sky130_fd_sc_hd__o2111ai_1
X_12476_ _03394_ net355 _03395_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__nand3_1
X_15264_ _06099_ _06093_ _06096_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__o21ai_2
X_11427_ _09526_ _02363_ _02356_ _02361_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__o211a_4
XPHY_EDGE_ROW_20_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14215_ _05037_ _05117_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__nand2_1
XANTENNA_5 _00127_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15195_ net739 net641 VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__nand2_1
X_11358_ _02293_ _02159_ _02291_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a21oi_2
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14146_ _04846_ _04843_ _04845_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_74_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ term_low\[23\] net1350 VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__nand2_1
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11289_ net228 _02132_ _02226_ _02227_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__o211ai_2
X_18954_ _09769_ _09770_ _09844_ _09845_ VGND VGND VPWR VPWR _09846_ sky130_fd_sc_hd__a22o_1
X_14077_ net778 net650 VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__nand2_1
X_17905_ _08762_ _08763_ VGND VGND VPWR VPWR _08764_ sky130_fd_sc_hd__and2_1
XFILLER_79_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13028_ _03953_ _03954_ _03949_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a21o_1
X_18885_ net596 net1001 VGND VGND VPWR VPWR _09777_ sky130_fd_sc_hd__nand2_1
X_17836_ _08695_ _08692_ _08687_ _08696_ VGND VGND VPWR VPWR _08697_ sky130_fd_sc_hd__o211ai_1
XFILLER_66_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer17 net812 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_89_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17767_ net960 net484 VGND VGND VPWR VPWR _08629_ sky130_fd_sc_hd__nand2_2
Xrebuffer28 net824 VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd1_1
X_14979_ _05757_ _05756_ _05754_ _05874_ _05873_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__o2111ai_4
Xrebuffer39 net835 VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_35_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19506_ _00586_ _00587_ _00692_ _00695_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__o22ai_2
X_16718_ _07450_ _07565_ _07564_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__a21boi_4
X_17698_ _08557_ _08559_ VGND VGND VPWR VPWR _08561_ sky130_fd_sc_hd__nor2_1
XFILLER_62_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16649_ _07376_ _07383_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__nand2_1
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19437_ _00616_ _00620_ _00619_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__a21o_1
XFILLER_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19368_ _05044_ _06521_ _10080_ _10106_ _10108_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__o2111ai_1
XFILLER_22_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18319_ _09140_ _09141_ _09163_ VGND VGND VPWR VPWR _09168_ sky130_fd_sc_hd__o21ai_1
Xrebuffer107 net903 VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer118 b_l\[10\] VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__buf_6
X_19299_ _00467_ _00469_ _00470_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__a21bo_1
Xrebuffer129 net765 VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd1_1
Xhold500 mid_sum\[23\] VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 mid_sum\[0\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 mid_sum\[32\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 p_lh\[31\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap252 _09225_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_1
X_20212_ _01350_ _01453_ _01454_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__a21oi_4
Xhold533 p_ll\[26\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 term_high\[60\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 p_lh\[0\] VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap263 _05741_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_6
Xmax_cap285 _05632_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_2
X_20143_ _01358_ _01380_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__xnor2_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20074_ _01299_ _01302_ _01304_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10660_ _01701_ _01702_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10591_ net793 net1325 VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__and2_1
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12330_ net906 net647 net511 net508 VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__nand4_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ _03183_ _03189_ _03190_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__nand3_2
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11212_ net691 net517 VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__and2_1
XFILLER_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14000_ _04746_ _04890_ _04899_ _04901_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__o22ai_4
X_12192_ _03006_ _03009_ _03010_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__a21o_1
X_11143_ _02081_ _02083_ _02078_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__a21oi_2
Xoutput75 net75 VGND VGND VPWR VPWR p[18] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput97 net97 VGND VGND VPWR VPWR p[38] sky130_fd_sc_hd__buf_2
X_15951_ _06824_ net262 VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__nand2_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11074_ net702 net517 VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__and2_1
Xoutput86 net86 VGND VGND VPWR VPWR p[28] sky130_fd_sc_hd__buf_2
X_15882_ _06757_ _06758_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__nand2_2
XFILLER_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18670_ _09345_ _09344_ _09342_ _09337_ VGND VGND VPWR VPWR _09551_ sky130_fd_sc_hd__o2bb2ai_2
X_14902_ _05796_ _05799_ _05800_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__a21oi_2
XFILLER_91_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17621_ _08484_ net476 net581 _08483_ VGND VGND VPWR VPWR _08485_ sky130_fd_sc_hd__and4_1
X_14833_ _05585_ _05732_ _05731_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_19_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11976_ _02908_ _02891_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__nand2_1
X_17552_ _08316_ _08325_ _08313_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__o21a_1
XFILLER_63_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14764_ _05263_ _05662_ _05664_ _05660_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__o211ai_1
X_10927_ _01873_ _01874_ _01867_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__a21bo_1
X_16503_ _07373_ _07374_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__nand2_1
X_17483_ _08346_ _08347_ _08342_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__a21oi_2
XFILLER_72_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13715_ _04604_ _04606_ _04614_ _04615_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__o2bb2ai_1
X_14695_ _05592_ _05595_ _05591_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__nand3_4
X_16434_ _07186_ _07307_ net797 VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__a21oi_1
XFILLER_71_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19222_ _10116_ net206 _10008_ VGND VGND VPWR VPWR _10120_ sky130_fd_sc_hd__a21o_1
XFILLER_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13646_ net741 net734 VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__nand2_8
X_10858_ net793 net1280 VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__and2_1
X_16365_ _06440_ _07234_ net561 net541 _07233_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__o2111ai_1
X_10789_ _01811_ _01812_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__nand2_1
X_13577_ _04431_ _04399_ _04430_ net1134 _04453_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__a32oi_4
XFILLER_31_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19153_ net562 net809 net776 net556 VGND VGND VPWR VPWR _10045_ sky130_fd_sc_hd__nand4_4
X_16296_ _07167_ _07169_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__nor2_1
X_18104_ _08894_ _08950_ _08952_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__a21boi_1
X_12528_ net292 _03453_ _03456_ _03418_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__o211ai_1
X_15316_ _06208_ _06209_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__nand2_1
X_19084_ _09970_ _09966_ _09906_ VGND VGND VPWR VPWR _09975_ sky130_fd_sc_hd__a21o_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12459_ _03387_ _03389_ _03383_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__a21o_1
X_18035_ _08882_ _08883_ _08857_ VGND VGND VPWR VPWR _08885_ sky130_fd_sc_hd__a21boi_2
X_15247_ _06081_ _06137_ _06138_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__nand3_1
XFILLER_125_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15178_ _05884_ _05985_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__nor2_2
XFILLER_99_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14129_ _05004_ _05030_ _05006_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__a21boi_1
X_19986_ _01208_ _01210_ net580 net721 VGND VGND VPWR VPWR _01212_ sky130_fd_sc_hd__and4_1
XFILLER_113_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18937_ _09806_ net446 _09804_ _09824_ _09826_ VGND VGND VPWR VPWR _09829_ sky130_fd_sc_hd__o2111ai_1
XFILLER_140_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18868_ _09605_ _09616_ _09755_ _09757_ VGND VGND VPWR VPWR _09760_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_38_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17819_ _08677_ _08678_ VGND VGND VPWR VPWR _08680_ sky130_fd_sc_hd__nand2_1
X_18799_ _09678_ _09689_ _09691_ VGND VGND VPWR VPWR _09692_ sky130_fd_sc_hd__nand3b_2
XFILLER_54_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20761_ clknet_leaf_53_clk _00401_ VGND VGND VPWR VPWR p_ll\[31\] sky130_fd_sc_hd__dfxtp_1
X_20692_ clknet_leaf_3_clk _00332_ VGND VGND VPWR VPWR p_hl\[26\] sky130_fd_sc_hd__dfxtp_2
XFILLER_10_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold374 p_hh_pipe\[6\] VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 p_hh\[2\] VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold396 p_ll_pipe\[2\] VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 p_ll\[22\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20126_ _01294_ _01360_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__nand2_1
X_20057_ _01205_ _01283_ net574 net721 _01286_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_146_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11830_ _02763_ _02765_ net712 net475 VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__and4_1
X_11761_ _02695_ _02696_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__or2_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_10712_ _01745_ _01746_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__nor2_1
X_13500_ _04348_ _04350_ _04352_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__o21ai_1
X_11692_ net664 net658 net526 net1059 VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__nand4_2
X_14480_ _05191_ _05194_ _05223_ _05381_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__o211ai_4
X_10643_ _01686_ _01687_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__nor2_1
X_13431_ _04339_ _04340_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_24_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16150_ net972 net1032 VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__nand2_1
XFILLER_139_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13362_ net766 net701 net693 net772 VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__a22o_1
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10574_ _09690_ net1338 VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__and2_1
X_16081_ net620 net502 VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__nand2_1
X_12313_ _03241_ _03244_ _03246_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__o21ai_4
XFILLER_6_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15101_ _05918_ _05960_ _05961_ _05915_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__a31o_1
XFILLER_142_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13293_ _04205_ _04157_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15032_ _05926_ _05927_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nand2_1
XFILLER_135_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12244_ _03041_ _03175_ a_h\[3\] net475 _03176_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__o2111a_1
XFILLER_107_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12175_ _03104_ _03106_ net226 _02940_ VGND VGND VPWR VPWR _03110_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_71_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19840_ _00895_ _01046_ _01049_ _01051_ VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__nand4_2
XFILLER_122_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11126_ net697 net517 _02066_ _02068_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__a22o_1
XFILLER_3_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19771_ net894 net556 VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__and2_1
X_16983_ _07593_ net477 net843 _07594_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__a31o_1
XFILLER_110_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18722_ _04555_ _06521_ VGND VGND VPWR VPWR _09607_ sky130_fd_sc_hd__nor2_1
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15934_ _06806_ _06811_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__nand2_1
X_11057_ _01961_ _02000_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__nand2_1
XFILLER_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15865_ a_l\[0\] net496 VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__nand2_1
X_18653_ _09405_ _09409_ _09407_ VGND VGND VPWR VPWR _09532_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_86_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17604_ _08415_ _08417_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__nand2_1
X_18584_ _09452_ net759 net597 VGND VGND VPWR VPWR _09456_ sky130_fd_sc_hd__nand3_1
X_14816_ net740 net663 VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__nand2_1
X_15796_ _06600_ _06607_ _06603_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_103_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17535_ _08399_ net488 a_l\[11\] VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__nand3_1
X_11959_ net644 net535 VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__nand2_1
X_14747_ _05546_ _05548_ _05643_ _05645_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__a22o_1
X_17466_ _08179_ _08190_ _08329_ _08331_ VGND VGND VPWR VPWR _08332_ sky130_fd_sc_hd__o211ai_1
X_14678_ _05573_ _05575_ _05569_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__a21o_1
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16417_ _07285_ _07286_ _07222_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__a21o_1
X_17397_ _08165_ _08262_ _08263_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__nand3_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13629_ _04535_ _04516_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_43_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19205_ _10092_ _10095_ _10079_ _10081_ _10098_ VGND VGND VPWR VPWR _10102_ sky130_fd_sc_hd__o221ai_4
XFILLER_146_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16348_ _07218_ _07220_ VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__nand2_1
X_19136_ _10024_ _10023_ _10011_ VGND VGND VPWR VPWR _10027_ sky130_fd_sc_hd__nand3_4
XFILLER_146_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16279_ _07152_ _07153_ _07089_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__a21oi_2
X_19067_ _09926_ _09954_ _09955_ VGND VGND VPWR VPWR _09958_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_113_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18018_ net459 _06521_ _08837_ _08840_ VGND VGND VPWR VPWR _08868_ sky130_fd_sc_hd__o22a_1
XFILLER_141_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19969_ _01143_ _01149_ _01190_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__and3_2
XFILLER_83_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20744_ clknet_leaf_42_clk _00384_ VGND VGND VPWR VPWR p_ll\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20675_ clknet_leaf_55_clk _00315_ VGND VGND VPWR VPWR p_hl\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire518 b_h\[5\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_21_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10290_ term_low\[20\] term_mid\[20\] VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__xnor2_1
XFILLER_12_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20109_ _01343_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__nand2b_1
X_13980_ net762 net670 _04877_ _04879_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a22o_1
X_12931_ _03802_ _03803_ _03857_ net175 VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__nand4_1
X_15650_ _06522_ _06524_ _09210_ _09581_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_100_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12862_ _03600_ _03702_ _03703_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__a21boi_4
X_11813_ _02745_ _02746_ _02730_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__a21o_1
X_14601_ _05463_ _05464_ _05499_ _05501_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_29_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ net631 net515 VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__nand2_1
X_12793_ net680 net474 _03719_ _03720_ VGND VGND VPWR VPWR _03722_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11744_ net951 _02679_ _02680_ _02467_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__o2bb2ai_1
X_17320_ _08177_ net341 _08183_ _08185_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14532_ _05428_ _05430_ _05431_ _05305_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__o2bb2ai_2
X_17251_ _08100_ net450 _08098_ _08116_ VGND VGND VPWR VPWR _08119_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ net854 net645 VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__nand2_8
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14463_ _05362_ _05363_ _05219_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__a21oi_2
XFILLER_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16202_ _09166_ _09657_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__nor2_1
X_17182_ _07812_ _07906_ _08045_ VGND VGND VPWR VPWR _08050_ sky130_fd_sc_hd__and3_1
X_10626_ p_hl\[0\] net1326 net797 VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__a21oi_1
X_13414_ _04271_ _04272_ _04273_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_40_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16133_ _06990_ _06994_ _07006_ _07008_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__nand4_1
X_14394_ _05170_ _05293_ _05292_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__nand4_4
X_10557_ net793 net1203 VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__and2_1
XFILLER_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13345_ _04215_ _04245_ _04247_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__o21ai_1
X_10488_ _01645_ term_high\[49\] net1345 VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__a21oi_1
X_16064_ _06937_ _06938_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__nand2_1
X_13276_ _04161_ _04165_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__nor2_1
Xrebuffer290 net792 VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12227_ _03004_ _03022_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__o21a_1
X_15015_ _05798_ _05803_ _05909_ _05910_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__o211ai_2
X_19823_ _01033_ _01029_ _01032_ _01004_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__o211ai_4
XFILLER_123_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12158_ _02852_ _03091_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__and3_1
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11109_ _01997_ _02047_ _02046_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__nand3_4
X_16966_ _07832_ _07805_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__nand2_2
X_12089_ _03002_ _03003_ _03016_ _03017_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__nand4_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19754_ _00960_ _00860_ _00959_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__nand3_1
X_15917_ net1127 net512 net505 net624 VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__a22oi_1
X_18705_ net153 _09312_ _09436_ _09313_ VGND VGND VPWR VPWR _09589_ sky130_fd_sc_hd__a22oi_2
X_19685_ _00747_ _00754_ _00882_ _00884_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__o22ai_4
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16897_ _07743_ _07745_ _07760_ _07762_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__a22o_1
X_18636_ _09506_ _09507_ _09494_ _09496_ VGND VGND VPWR VPWR _09513_ sky130_fd_sc_hd__o211ai_4
X_15848_ _06636_ _06641_ _06724_ _06725_ VGND VGND VPWR VPWR _06727_ sky130_fd_sc_hd__nand4_2
XFILLER_80_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15779_ net624 net512 VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__nand2_1
X_18567_ _09436_ _09437_ VGND VGND VPWR VPWR _09438_ sky130_fd_sc_hd__and2_1
X_17518_ _08382_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__inv_2
X_18498_ _04182_ _06867_ _09354_ VGND VGND VPWR VPWR _09363_ sky130_fd_sc_hd__o21ba_4
XFILLER_33_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17449_ _08308_ _08310_ _08304_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__a21o_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20460_ clknet_leaf_14_clk _00100_ VGND VGND VPWR VPWR term_high\[52\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_115_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20391_ clknet_leaf_37_clk _00031_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfxtp_1
X_19119_ _09253_ _09275_ net457 _09915_ VGND VGND VPWR VPWR _10009_ sky130_fd_sc_hd__o31a_1
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20727_ clknet_leaf_7_clk _00367_ VGND VGND VPWR VPWR p_lh\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20658_ clknet_leaf_12_clk _00298_ VGND VGND VPWR VPWR p_hh\[24\] sky130_fd_sc_hd__dfxtp_1
Xwire326 _02574_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
X_11460_ _09406_ _09613_ _02256_ _02397_ _02396_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__o221ai_2
XFILLER_109_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10411_ term_mid\[37\] term_high\[37\] term_mid\[36\] term_high\[36\] VGND VGND VPWR
+ VPWR _01582_ sky130_fd_sc_hd__o211a_1
X_11391_ _02331_ _02330_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__nand2_4
XFILLER_137_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20589_ clknet_leaf_14_clk _00229_ VGND VGND VPWR VPWR p_hh_pipe\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_99_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13130_ _04013_ _04050_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__nand2_1
X_10342_ _00891_ _00956_ _00967_ _01042_ VGND VGND VPWR VPWR _01139_ sky130_fd_sc_hd__or4b_1
XFILLER_140_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13061_ _03984_ _03976_ _03983_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__nand3_1
X_12012_ net247 _02942_ _02945_ _02937_ _02936_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__o2111ai_2
X_10273_ term_low\[18\] term_mid\[18\] VGND VGND VPWR VPWR _10126_ sky130_fd_sc_hd__nor2_1
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16820_ _07684_ _07687_ _07664_ net278 VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__o211ai_2
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16751_ _07478_ _07467_ _07469_ VGND VGND VPWR VPWR _07622_ sky130_fd_sc_hd__o21a_1
XFILLER_93_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone216 net564 VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__clkbuf_16
X_15702_ _06538_ _06578_ _06579_ _06580_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__or4_4
XFILLER_46_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13963_ _04862_ _04867_ _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__o21ai_2
X_16682_ _07491_ _07551_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__nand2_1
X_12914_ _03815_ _03817_ _03836_ _03837_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__a22o_1
X_13894_ _04797_ _04798_ _04667_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nand3_1
X_19470_ _00455_ _00653_ _00656_ _00652_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__o211ai_2
X_15633_ _06474_ _06483_ _06484_ _06490_ _06472_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__a32o_1
XFILLER_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12845_ _03727_ _03772_ _03773_ VGND VGND VPWR VPWR _03774_ sky130_fd_sc_hd__nand3_2
X_18421_ _09274_ _09276_ _09269_ VGND VGND VPWR VPWR _09279_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12776_ _03600_ _03609_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__nand2_1
X_15564_ _06446_ net423 _06444_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__nand3_2
X_18352_ _09200_ _09198_ _09111_ VGND VGND VPWR VPWR _09204_ sky130_fd_sc_hd__nand3_2
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11727_ _02647_ _02644_ _02660_ _02661_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__o2bb2ai_4
X_17303_ _02338_ _07234_ VGND VGND VPWR VPWR _08170_ sky130_fd_sc_hd__nor2_1
X_14515_ _02613_ _04182_ _05270_ _05273_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__o22a_4
XFILLER_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18283_ net457 _06441_ _09030_ _09124_ _09125_ VGND VGND VPWR VPWR _09129_ sky130_fd_sc_hd__o2111ai_1
X_15495_ _06365_ _06345_ _06384_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__o21ai_1
XFILLER_14_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11658_ _02586_ _02585_ _02592_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__a21o_1
X_17234_ _07951_ _07954_ _02338_ _06985_ VGND VGND VPWR VPWR _08102_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_80_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14446_ _05348_ net690 net730 VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__nand3_1
X_11589_ _09417_ _09613_ _02526_ _02527_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__o211ai_2
X_17165_ _07967_ _07969_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__nor2_1
X_10609_ net794 net1220 VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__and2_1
X_14377_ net761 net655 _05274_ _05275_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__a22o_1
XFILLER_142_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16116_ _06983_ _06986_ _09286_ _09581_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__o2bb2ai_1
Xmax_cap615 net616 VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__buf_12
Xmax_cap604 net606 VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__buf_8
X_13328_ _04239_ _04240_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__nand2_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17096_ _07964_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__inv_2
Xmax_cap637 net638 VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__buf_12
Xmax_cap659 net661 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_8
X_16047_ _06890_ _06915_ _06913_ _06894_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__o211ai_2
XFILLER_124_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13259_ _04171_ _04172_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__nand3_2
XFILLER_97_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19806_ net1033 net567 net1013 net1079 VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__a22o_1
X_17998_ _08833_ _08847_ VGND VGND VPWR VPWR _08849_ sky130_fd_sc_hd__or2_1
X_19737_ _00939_ _00940_ _00941_ _00810_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__o2bb2ai_2
X_16949_ net558 net523 net516 net566 VGND VGND VPWR VPWR _07819_ sky130_fd_sc_hd__a22oi_4
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19668_ net893 net563 VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__nand2_1
XFILLER_80_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18619_ _09488_ _09477_ VGND VGND VPWR VPWR _09495_ sky130_fd_sc_hd__nand2_1
XFILLER_52_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19599_ net579 net738 VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_121_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20512_ clknet_leaf_35_clk _00152_ VGND VGND VPWR VPWR term_low\[7\] sky130_fd_sc_hd__dfxtp_1
X_20443_ clknet_leaf_28_clk _00083_ VGND VGND VPWR VPWR term_high\[35\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20374_ clknet_leaf_52_clk _00014_ VGND VGND VPWR VPWR b_l\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_133_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10960_ _01895_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__nor2_1
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10891_ net794 net1159 VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__and2_1
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12630_ _03548_ _03557_ _03549_ VGND VGND VPWR VPWR _03561_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_48_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12561_ _03357_ _03363_ _03377_ _03487_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__a22oi_1
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11512_ net708 net487 VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__and2_1
X_12492_ net633 b_h\[4\] net518 net1049 VGND VGND VPWR VPWR _03424_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _06167_ _06169_ _06159_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__o21bai_2
X_14300_ net740 net685 VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__nand2_1
Xwire134 _00073_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
X_11443_ _02370_ _02372_ _02382_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__a21o_1
Xwire156 _06207_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14231_ _05121_ _05131_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__nand2_1
Xwire178 _02678_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__buf_1
Xwire167 _01471_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__buf_2
X_14162_ net350 _05066_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__nand2_1
X_11374_ _02184_ _02250_ _02313_ _02314_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__o211ai_4
X_13113_ _04035_ _03953_ _04037_ VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__a21boi_2
XFILLER_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18970_ _09860_ _09861_ VGND VGND VPWR VPWR _09862_ sky130_fd_sc_hd__or2_1
X_10325_ term_low\[26\] term_mid\[26\] VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__and2_1
X_14093_ _04990_ _04993_ _04997_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__o21ai_1
X_10256_ _09690_ net1186 VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__and2_1
X_17921_ _08722_ _08723_ _08750_ _08753_ VGND VGND VPWR VPWR _08779_ sky130_fd_sc_hd__a31o_1
XFILLER_79_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _03904_ _03905_ _03965_ _03967_ _03910_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__o221ai_4
XFILLER_121_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17852_ _08619_ net137 _08669_ _08614_ VGND VGND VPWR VPWR _08713_ sky130_fd_sc_hd__o211ai_1
XFILLER_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16803_ _07670_ _07672_ net590 net503 VGND VGND VPWR VPWR _07674_ sky130_fd_sc_hd__and4_1
X_10187_ net926 VGND VGND VPWR VPWR _09220_ sky130_fd_sc_hd__inv_12
XFILLER_94_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17783_ _08644_ _08642_ _08641_ VGND VGND VPWR VPWR _08645_ sky130_fd_sc_hd__nand3_1
X_14995_ _05874_ _05876_ _05873_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__a21boi_4
X_16734_ net950 net496 VGND VGND VPWR VPWR _07605_ sky130_fd_sc_hd__nand2_1
X_19522_ _10004_ _00711_ _10002_ _00713_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__a31o_1
X_13946_ _04845_ _04846_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__nand2_1
X_16665_ _07533_ _07535_ _07521_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__and3_1
X_19453_ b_l\[3\] net811 net552 net548 VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__nand4_4
X_15616_ _06493_ _06496_ _06431_ _06432_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__o2bb2ai_1
X_18404_ _09243_ _09247_ _09259_ VGND VGND VPWR VPWR _09260_ sky130_fd_sc_hd__nand3_1
XFILLER_50_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13877_ net741 net734 net703 net701 VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__nand4_4
X_16596_ _07463_ _07464_ _07466_ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__nand3_1
X_12828_ _03754_ _03756_ VGND VGND VPWR VPWR _03757_ sky130_fd_sc_hd__nand2_1
X_19384_ _00561_ _00562_ _00563_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _06404_ _06418_ _06420_ _06421_ _06411_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__a32o_1
X_12759_ _03452_ _03531_ _03567_ _03687_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o22ai_2
X_18335_ _09169_ _09175_ _09180_ _09178_ VGND VGND VPWR VPWR _09185_ sky130_fd_sc_hd__o211ai_4
XFILLER_61_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18266_ _09089_ _09091_ net373 _09087_ VGND VGND VPWR VPWR _09112_ sky130_fd_sc_hd__a2bb2oi_1
X_15478_ _06314_ _06315_ _06349_ _06353_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_96_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17217_ _08073_ _08078_ _08081_ VGND VGND VPWR VPWR _08085_ sky130_fd_sc_hd__a21oi_1
X_14429_ _05330_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__nand2_2
X_18197_ _09041_ _09038_ _09039_ VGND VGND VPWR VPWR _09044_ sky130_fd_sc_hd__a21oi_1
XFILLER_116_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17148_ _08009_ _08011_ _08013_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap445 _00747_ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__buf_6
XFILLER_143_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap467 _01762_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
X_17079_ _07634_ _07789_ _07803_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__o21ai_2
Xmax_cap478 b_h\[14\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__buf_8
Xmax_cap456 _04608_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_2
XFILLER_112_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap489 net490 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_8
X_20090_ net580 b_l\[15\] VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__nand2_1
XFILLER_130_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_49_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_123_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20426_ clknet_leaf_14_clk net1346 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20357_ net794 net54 VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__and2_1
X_11090_ _01970_ _01998_ _02031_ _02032_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__o211ai_2
XFILLER_121_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20288_ _01532_ _01533_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11992_ _02918_ _02921_ _02861_ _02920_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__o211ai_4
XFILLER_91_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14780_ net745 net655 VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__nand2_1
X_13800_ net752 net683 VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__nand2_2
X_10943_ net691 net545 net538 net697 VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__a22oi_2
X_13731_ _04633_ _04636_ _04631_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__o21bai_2
XFILLER_16_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16450_ net928 net496 VGND VGND VPWR VPWR _07323_ sky130_fd_sc_hd__nand2_1
X_10874_ _09690_ net1172 VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__and2_1
X_13662_ _04568_ _04566_ _04569_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__a21o_1
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16381_ _07242_ _07249_ _07248_ _07240_ _07241_ VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__o2111ai_1
X_12613_ _09471_ _09646_ _03539_ _03541_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__o211ai_1
X_13593_ _04498_ _04499_ _04488_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__a21o_1
X_15401_ _06292_ _06293_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ _03470_ _03471_ _03474_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__a21oi_1
X_18120_ net781 net601 net594 net790 VGND VGND VPWR VPWR _08968_ sky130_fd_sc_hd__a22oi_1
XFILLER_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15332_ net719 net657 _06223_ _06224_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__a22o_1
XFILLER_129_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18051_ _08899_ VGND VGND VPWR VPWR _08900_ sky130_fd_sc_hd__inv_2
XFILLER_12_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17002_ _07868_ _07869_ _07871_ VGND VGND VPWR VPWR _07872_ sky130_fd_sc_hd__a21o_1
X_12475_ net355 _03394_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15263_ _06154_ _06156_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__nand2_1
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_6 _00296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11426_ _02361_ _02364_ _02356_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__a21o_1
X_14214_ _04968_ _05031_ net244 _05039_ _05081_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__a32oi_2
X_15194_ _05797_ net635 net745 VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__and3_2
X_11357_ _02295_ _02296_ _09428_ _09602_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o2bb2ai_1
X_14145_ _05048_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_91_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18953_ _09839_ _09772_ _09838_ VGND VGND VPWR VPWR _09845_ sky130_fd_sc_hd__nand3_2
XFILLER_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ _00676_ _00730_ _00698_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__o21ai_1
X_14076_ _04892_ _04898_ _04895_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__a21oi_1
X_11288_ net228 _02132_ _02226_ _02227_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__o211a_1
X_17904_ _09319_ _09679_ _08726_ VGND VGND VPWR VPWR _08763_ sky130_fd_sc_hd__or3b_1
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13027_ _03950_ _03952_ _03951_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__nand3_1
X_18884_ net1111 net747 VGND VGND VPWR VPWR _09776_ sky130_fd_sc_hd__nand2_1
X_10239_ net794 net63 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__and2_1
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17835_ _08691_ _08693_ _08688_ VGND VGND VPWR VPWR _08696_ sky130_fd_sc_hd__a21o_1
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer18 net812 VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__buf_2
X_17766_ _08596_ _08599_ VGND VGND VPWR VPWR _08628_ sky130_fd_sc_hd__and2_1
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16717_ _07450_ _07565_ _07560_ _07563_ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_89_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer29 net824 VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd1_1
X_14978_ net1147 _05874_ _05875_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__a21o_1
X_19505_ _00685_ _00694_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__nor2_4
XFILLER_90_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17697_ net1093 net476 _08552_ _08555_ VGND VGND VPWR VPWR _08560_ sky130_fd_sc_hd__a22o_1
X_13929_ _04774_ _04801_ _04803_ _04775_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__a31oi_1
XFILLER_34_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16648_ _07514_ _07518_ _07517_ VGND VGND VPWR VPWR _07520_ sky130_fd_sc_hd__o21a_1
XFILLER_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19436_ _09199_ _09362_ _00612_ _00613_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__o22a_1
X_16579_ _07348_ _07416_ _07414_ VGND VGND VPWR VPWR _07451_ sky130_fd_sc_hd__a21oi_2
X_19367_ _10077_ _10080_ _10105_ _10107_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_TAPCELL_ROW_33_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18318_ _09161_ _09162_ _09145_ VGND VGND VPWR VPWR _09167_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_100_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer108 b_h\[1\] VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer119 net915 VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd1_1
X_19298_ net1065 _00469_ _00470_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__a21boi_1
X_18249_ net187 _09094_ net207 VGND VGND VPWR VPWR _09096_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold501 mid_sum\[7\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 term_high\[53\] VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 term_high\[54\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap253 net254 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
Xhold512 mid_sum\[31\] VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
X_20211_ _01344_ _01401_ _01403_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__o21ai_2
XFILLER_104_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold567 _00178_ VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 p_lh\[30\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap275 _09416_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_1
Xmax_cap264 _04562_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__buf_1
X_20142_ _01378_ _01379_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__nand2_1
XFILLER_98_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20073_ _01297_ _01301_ _01304_ _01299_ VGND VGND VPWR VPWR _01306_ sky130_fd_sc_hd__o211ai_4
XFILLER_100_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10590_ net793 net1301 VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__and2_1
XFILLER_21_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12260_ _03192_ _03182_ _03191_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__nand3_2
X_20409_ clknet_leaf_29_clk _00049_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfxtp_1
X_12191_ _03037_ _03080_ _03034_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__a21oi_4
X_11211_ _02073_ _02091_ _02092_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__a21boi_4
X_11142_ _02083_ net534 net681 VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__nand3_1
XFILLER_1_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput76 net76 VGND VGND VPWR VPWR p[19] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput98 net98 VGND VGND VPWR VPWR p[39] sky130_fd_sc_hd__buf_2
X_15950_ _06745_ _06747_ _06824_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__o21ai_2
X_11073_ _02002_ _02010_ _02012_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__nand3_2
Xoutput87 net87 VGND VGND VPWR VPWR p[29] sky130_fd_sc_hd__buf_2
X_15881_ net595 net531 net527 net602 VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__a22oi_1
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14901_ net745 net649 VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__and2_1
X_17620_ _08480_ _08481_ VGND VGND VPWR VPWR _08484_ sky130_fd_sc_hd__nand2_1
X_14832_ _05712_ _05713_ _05726_ _05727_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__nand4_2
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _02890_ _02885_ _02889_ net323 _02907_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__o2111ai_4
XFILLER_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17551_ _08413_ _08415_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__nand2_1
XFILLER_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14763_ _05408_ _05533_ _05531_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__a21o_1
X_10926_ _01868_ _01870_ _01872_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__nand3_1
X_16502_ net561 net533 net529 net570 VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__a22oi_2
X_17482_ _08346_ _08342_ _08347_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__and3_1
X_13714_ _04599_ _04605_ _04618_ _04604_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__o211ai_1
X_14694_ _05458_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nand2_2
X_16433_ _07167_ _07169_ _07175_ _07304_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__o41a_1
X_10857_ net793 net1266 VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__and2_1
X_13645_ net741 net734 VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__and2_1
X_19221_ net206 _10116_ _10008_ VGND VGND VPWR VPWR _10119_ sky130_fd_sc_hd__a21oi_2
X_19152_ _09942_ _10042_ VGND VGND VPWR VPWR _10044_ sky130_fd_sc_hd__nand2_2
X_16364_ _07233_ _07235_ _09319_ _09581_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__o2bb2ai_1
X_10788_ _01794_ _01796_ _01803_ _01809_ _01802_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__a311oi_1
X_18103_ _08946_ _08948_ _08894_ _09690_ VGND VGND VPWR VPWR _08952_ sky130_fd_sc_hd__o31a_1
X_13576_ _04479_ _04387_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16295_ _07166_ net282 _07165_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__nand3_4
X_12527_ _03449_ _03454_ _03456_ net246 _03415_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__o2111ai_4
X_15315_ _06209_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__inv_2
X_19083_ _09906_ _09966_ _09970_ VGND VGND VPWR VPWR _09974_ sky130_fd_sc_hd__nand3_2
X_12458_ _03387_ _03389_ _03383_ VGND VGND VPWR VPWR _03390_ sky130_fd_sc_hd__a21oi_1
X_18034_ _08882_ _08883_ VGND VGND VPWR VPWR _08884_ sky130_fd_sc_hd__nand2_1
X_15246_ _06137_ _06138_ _06081_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__a21o_1
X_11409_ _02264_ _02265_ _02263_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__a21bo_1
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12389_ _03317_ net460 _03308_ _03316_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__o211a_1
X_15177_ _05982_ _05882_ _05983_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__a21o_1
X_19985_ _01210_ net721 net580 VGND VGND VPWR VPWR _01211_ sky130_fd_sc_hd__and3_1
X_14128_ _05000_ _05005_ _05032_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14059_ _04694_ _04829_ net142 _04824_ _04693_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__o32a_1
X_18936_ _09808_ _09824_ _09826_ VGND VGND VPWR VPWR _09828_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18867_ _09605_ _09616_ _09755_ _09757_ VGND VGND VPWR VPWR _09759_ sky130_fd_sc_hd__o22a_1
X_17818_ net962 net555 net486 net999 VGND VGND VPWR VPWR _08679_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_38_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18798_ _09684_ _09685_ _09680_ VGND VGND VPWR VPWR _09691_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_38_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17749_ _08609_ _08610_ _08611_ VGND VGND VPWR VPWR _08612_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20760_ clknet_leaf_53_clk _00400_ VGND VGND VPWR VPWR p_ll\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19419_ net588 net579 net744 net738 _00595_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__a41o_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20691_ clknet_leaf_3_clk _00331_ VGND VGND VPWR VPWR p_hl\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold364 term_low\[8\] VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold375 p_ll\[2\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 p_ll\[1\] VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold397 term_low\[11\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
X_20125_ net731 net549 VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__nand2_1
X_20056_ _01286_ net721 net574 _01285_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__and4_1
XFILLER_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _02695_ _02696_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__nor2_1
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ _01742_ _01743_ _01744_ net796 VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__a31o_1
XFILLER_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11691_ net664 net658 net526 net1059 VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__and4_1
X_10642_ p_hl\[3\] p_lh\[3\] VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__and2_1
X_13430_ net766 net693 net986 net923 VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_24_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ net766 net701 net693 net923 VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__a22oi_1
X_10573_ _09690_ net1336 VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__and2_1
X_12312_ _02967_ _03099_ _03100_ _03106_ _03109_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__a32o_1
XFILLER_127_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16080_ net607 _06879_ net515 _06881_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__a31o_4
X_13292_ _04204_ _04205_ _04157_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer9 _05574_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd1_1
X_15100_ _05994_ _05995_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__nand2_1
X_12243_ net687 net483 _03043_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_58_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15031_ net733 net657 net651 net739 VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__a22oi_2
X_12174_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__inv_2
XFILLER_122_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_71_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11125_ net691 net1078 net525 net519 VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__nand4_2
X_16982_ _07695_ _07733_ _07845_ _07847_ VGND VGND VPWR VPWR _07852_ sky130_fd_sc_hd__o22ai_2
XFILLER_68_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19770_ _00867_ _00953_ _00954_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__a21oi_2
X_15933_ _06790_ _06807_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__nand2_1
X_11056_ _01959_ _01963_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__nand2_1
X_18721_ _09603_ _09604_ VGND VGND VPWR VPWR _09606_ sky130_fd_sc_hd__nand2_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15864_ _06582_ _06721_ _06719_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__a21oi_4
X_18652_ _09405_ _09409_ _09407_ VGND VGND VPWR VPWR _09531_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15795_ net382 _06615_ _06614_ net1007 VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__a2bb2oi_2
X_17603_ net581 net1093 _02588_ _08388_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__a31o_1
X_18583_ _09453_ net1001 net606 VGND VGND VPWR VPWR _09455_ sky130_fd_sc_hd__nand3_1
X_14815_ net730 net865 VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__nand2_1
XFILLER_91_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17534_ net565 net560 net500 net494 VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__nand4_2
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14746_ _05551_ _05641_ _05549_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__a21o_1
X_11958_ _09515_ _09592_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__nor2_1
X_10909_ _09526_ _09581_ _01855_ _01858_ net795 VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__o311a_1
X_11889_ _02701_ _02715_ _02714_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o21ai_1
X_17465_ _08316_ _08325_ _08327_ _08324_ VGND VGND VPWR VPWR _08331_ sky130_fd_sc_hd__o211ai_4
X_19204_ _10092_ _10095_ _10098_ _10082_ _10080_ VGND VGND VPWR VPWR _10101_ sky130_fd_sc_hd__o2111ai_2
X_14677_ _09264_ _09482_ _05573_ _05575_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__o211ai_2
X_16416_ _07222_ _07285_ _07286_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__nand3_1
X_17396_ _08240_ _08244_ _08257_ _08258_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__o2bb2ai_1
X_13628_ _04514_ _04509_ net1050 _04530_ _04534_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_43_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16347_ _07212_ _07219_ _07217_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__a21oi_2
X_13559_ _04396_ net1133 _04463_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nand3_1
X_19135_ _10012_ _10021_ _10022_ VGND VGND VPWR VPWR _10026_ sky130_fd_sc_hd__nand3_1
XFILLER_146_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19066_ _09950_ _09952_ _09925_ VGND VGND VPWR VPWR _09957_ sky130_fd_sc_hd__a21oi_2
XFILLER_146_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16278_ _07123_ _07126_ _07128_ _07149_ VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__o211ai_4
X_18017_ _08837_ _08840_ _08839_ VGND VGND VPWR VPWR _08867_ sky130_fd_sc_hd__o21ai_2
XFILLER_126_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15229_ _06118_ _06119_ _06120_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_113_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19968_ _01127_ _01131_ _01142_ _01191_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__o211ai_4
X_19899_ _01017_ _01018_ _01022_ _01016_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__a22oi_1
X_18919_ net780 net1084 VGND VGND VPWR VPWR _09811_ sky130_fd_sc_hd__nand2_1
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20743_ clknet_leaf_42_clk _00383_ VGND VGND VPWR VPWR p_ll\[13\] sky130_fd_sc_hd__dfxtp_1
X_20674_ clknet_leaf_5_clk _00314_ VGND VGND VPWR VPWR p_hl\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20108_ _01262_ _01277_ _01340_ _01341_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__nand4_2
X_12930_ _03855_ _03856_ _03734_ _03771_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_46_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20039_ net203 _01264_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__nor2_2
X_12861_ _03786_ _03789_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__and2_1
XFILLER_74_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11812_ _02747_ _02730_ VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__nand2_1
X_14600_ _05465_ _05497_ _05498_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_29_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _06435_ _06448_ _06447_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__o21ai_1
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12792_ _03719_ _03720_ _03716_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _02468_ net402 _02243_ _02469_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__a31o_1
X_14531_ _05424_ _05429_ _05432_ _05428_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__o211ai_2
XFILLER_14_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11674_ _02609_ _02610_ VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__nand2_2
X_17250_ _08117_ _08101_ VGND VGND VPWR VPWR _08118_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _05220_ _05362_ _05363_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__and3_1
X_16201_ _07071_ _07067_ _07065_ _07070_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__o211ai_2
X_17181_ _07642_ _07811_ _08043_ _08044_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_81_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _01860_ _04260_ net714 net748 _04322_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_40_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ net794 net1282 VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16132_ _06998_ _07001_ _06995_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__a21o_1
X_14393_ _05155_ _05168_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__nand2_1
X_10556_ net793 net1233 VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__and2_1
XFILLER_128_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13344_ _04209_ _04210_ _04255_ _04256_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__o31a_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10487_ term_high\[49\] _01645_ _01646_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__o21a_1
XFILLER_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16063_ _06934_ _06936_ _06743_ _06744_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_115_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13275_ _09177_ _04187_ _04186_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__o21ai_1
Xrebuffer291 net792 VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer280 net1076 VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd1_1
X_12226_ _03157_ _03159_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__nand2_1
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15014_ _05905_ _05909_ _05910_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__and3_1
X_12157_ _02825_ _02847_ _02848_ _02854_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__a31o_1
XFILLER_69_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19822_ _01034_ _01003_ _01035_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__nand3_4
X_11108_ _01996_ net249 _02050_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__nand3_4
XFILLER_69_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16965_ _07800_ _07801_ _07830_ _07831_ VGND VGND VPWR VPWR _07835_ sky130_fd_sc_hd__o211ai_2
X_12088_ _03012_ _03014_ _03002_ VGND VGND VPWR VPWR _03023_ sky130_fd_sc_hd__o21ai_1
X_19753_ _00957_ _00958_ _00861_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__a21oi_1
X_15916_ net617 net512 VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__nand2_2
X_11039_ net466 _01912_ net712 net1018 VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__and4b_2
X_16896_ _07737_ _07764_ _07765_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__nand3_2
X_18704_ _09586_ _09580_ _09585_ VGND VGND VPWR VPWR _09588_ sky130_fd_sc_hd__a21o_1
X_19684_ _09319_ _09340_ net457 _00743_ net445 VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__o32a_4
X_15847_ _06722_ _06723_ _06653_ VGND VGND VPWR VPWR _06726_ sky130_fd_sc_hd__a21oi_1
X_18635_ _09510_ _09474_ _09509_ VGND VGND VPWR VPWR _09512_ sky130_fd_sc_hd__nand3_4
XFILLER_91_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15778_ net632 net502 VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__nand2_1
X_18566_ _09432_ _09434_ _09435_ VGND VGND VPWR VPWR _09437_ sky130_fd_sc_hd__nand3_4
X_17517_ _08379_ _08380_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__or2_2
X_18497_ net764 net1111 _09357_ _09360_ VGND VGND VPWR VPWR _09361_ sky130_fd_sc_hd__a22oi_2
X_14729_ _05608_ _05625_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__nand2_1
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17448_ _08305_ _08306_ _08304_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__o21ai_2
XFILLER_60_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17379_ _07962_ _08087_ _08123_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__o21ai_1
X_19118_ _09969_ _09967_ _09966_ _09906_ VGND VGND VPWR VPWR _10008_ sky130_fd_sc_hd__a22oi_4
XFILLER_145_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20390_ clknet_leaf_41_clk _00030_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19049_ net919 net568 net1084 net776 VGND VGND VPWR VPWR _09940_ sky130_fd_sc_hd__a22oi_2
XFILLER_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20726_ clknet_leaf_7_clk _00366_ VGND VGND VPWR VPWR p_lh\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10410_ _01570_ _01575_ _01565_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__and3_1
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire327 _02388_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_2
X_20657_ clknet_leaf_11_clk _00297_ VGND VGND VPWR VPWR p_hh\[23\] sky130_fd_sc_hd__dfxtp_1
Xwire316 _05076_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_1
X_11390_ net200 _02325_ _02230_ _02235_ net179 VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__o221ai_4
X_20588_ clknet_leaf_14_clk _00228_ VGND VGND VPWR VPWR p_hh_pipe\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10341_ term_low\[27\] term_mid\[27\] _01117_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a21o_1
X_10272_ _10018_ _10072_ _10061_ VGND VGND VPWR VPWR _10115_ sky130_fd_sc_hd__o21ai_2
X_13060_ _03983_ _03984_ _03976_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__a21o_1
XFILLER_2_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12011_ _02936_ _02937_ _02943_ _02944_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_105_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_131_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16750_ _07592_ _07618_ _07619_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__nand3b_4
Xclone239 net638 VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__clkbuf_16
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13962_ _04865_ _04866_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__nand2_1
X_15701_ _06540_ _06535_ _06578_ _06579_ _06538_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__a2111oi_4
X_12913_ _03815_ _03817_ _03836_ _03837_ VGND VGND VPWR VPWR _03841_ sky130_fd_sc_hd__nand4_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16681_ _07507_ _07508_ _07546_ _07547_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__nand4_1
X_18420_ _09274_ _09276_ _09270_ VGND VGND VPWR VPWR _09278_ sky130_fd_sc_hd__a21o_1
XFILLER_62_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13893_ _04797_ _04798_ _04667_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__and3_4
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15632_ _06474_ _06483_ _06484_ _06490_ _06472_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__a32oi_4
XFILLER_104_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _03734_ _03766_ _03767_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__nand3_2
XFILLER_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15563_ _06439_ _06442_ _06437_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__a21o_1
X_12775_ _03702_ _03703_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__nand2_1
X_18351_ _09186_ _09195_ _09112_ VGND VGND VPWR VPWR _09203_ sky130_fd_sc_hd__a21oi_1
X_11726_ _02662_ _02663_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__nand2_1
X_17302_ net569 net498 net493 net573 VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__a22oi_2
X_18282_ _09113_ _09124_ _09125_ VGND VGND VPWR VPWR _09128_ sky130_fd_sc_hd__nand3_2
X_14514_ _05270_ _05273_ _05275_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__o21ai_2
XFILLER_30_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_140_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17233_ net450 _08100_ _08098_ VGND VGND VPWR VPWR _08101_ sky130_fd_sc_hd__o21ai_2
X_15494_ _06382_ _06383_ VGND VGND VPWR VPWR _06384_ sky130_fd_sc_hd__nand2b_1
X_11657_ _02585_ _02586_ _02593_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__nand3_1
X_14445_ net740 net736 net685 net677 VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nand4_2
X_11588_ _02397_ net510 net681 VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__nand3_1
X_17164_ net612 net472 VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__nand2_1
X_10608_ net794 net1252 VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _05274_ _05275_ _05270_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__a21o_1
X_10539_ net793 net1226 VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__and2_1
XFILLER_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap616 net617 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__buf_12
X_16115_ _06983_ _06986_ net572 net541 VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__nand4_1
Xmax_cap605 net608 VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__buf_6
Xmax_cap627 net628 VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__buf_12
X_17095_ _07959_ _07961_ _07949_ VGND VGND VPWR VPWR _07964_ sky130_fd_sc_hd__nand3_4
X_13327_ _04238_ net710 net763 _04236_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__nand4_1
X_16046_ _06894_ _06913_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__nand2_2
Xmax_cap638 net641 VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__buf_12
Xmax_cap649 net650 VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__buf_8
XFILLER_6_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13258_ _04144_ _04151_ _04152_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__o21ai_1
X_12209_ _03138_ _03139_ _03140_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__nand3_1
X_13189_ _04082_ _04084_ _04105_ _04106_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__and4_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17997_ _08847_ _08833_ VGND VGND VPWR VPWR _08848_ sky130_fd_sc_hd__nand2_1
XFILLER_69_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19805_ b_l\[9\] net563 VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__nand2_1
X_16948_ _07815_ _07817_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__nand2_1
X_19736_ _00939_ _00940_ _00942_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_125_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16879_ net600 net488 VGND VGND VPWR VPWR _07749_ sky130_fd_sc_hd__nand2_1
X_19667_ _00772_ _00776_ _00831_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__o21ai_2
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18618_ _09372_ _09476_ _09491_ _09492_ VGND VGND VPWR VPWR _09494_ sky130_fd_sc_hd__o211ai_2
X_19598_ _00595_ _00601_ _00598_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__a21o_1
XFILLER_25_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18549_ _09412_ _09413_ _09415_ VGND VGND VPWR VPWR _09419_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20511_ clknet_leaf_32_clk _00151_ VGND VGND VPWR VPWR term_low\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20442_ clknet_leaf_28_clk _00082_ VGND VGND VPWR VPWR term_high\[34\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20373_ clknet_leaf_52_clk _00013_ VGND VGND VPWR VPWR b_l\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10890_ net794 net1208 VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__and2_1
XFILLER_70_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12560_ _03488_ _03489_ _03490_ VGND VGND VPWR VPWR _03492_ sky130_fd_sc_hd__a21o_1
X_11511_ _09624_ _09635_ _01860_ _02341_ _02342_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__o32a_1
X_12491_ net633 b_h\[4\] net518 net1049 VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__a22oi_1
X_20709_ clknet_leaf_40_clk _00349_ VGND VGND VPWR VPWR p_lh\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire135 _00348_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
X_11442_ _02379_ _02381_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__nand2_1
Xwire157 _04954_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14230_ _05121_ _05129_ _05130_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nand3b_4
Xwire179 _02324_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__buf_1
X_11373_ _02268_ _02269_ _02309_ _02310_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__a22o_1
X_14161_ _05059_ _05060_ _05051_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__nand3_1
X_13112_ _03993_ _03948_ _03995_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__o21a_1
X_10324_ _00913_ _00924_ _00935_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__a21oi_1
X_14092_ _04996_ _04980_ _04995_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nand3_2
X_10255_ _09690_ net1161 VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__and2_1
X_17920_ _08770_ _08777_ _08778_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_76_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _03902_ _03907_ _03906_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__o21ai_2
X_17851_ _08711_ VGND VGND VPWR VPWR _08712_ sky130_fd_sc_hd__inv_2
X_10186_ net606 VGND VGND VPWR VPWR _09210_ sky130_fd_sc_hd__inv_8
X_16802_ _07670_ _07672_ _09253_ _09613_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__o2bb2ai_1
X_17782_ _08562_ _08574_ _08576_ VGND VGND VPWR VPWR _08644_ sky130_fd_sc_hd__o21ai_2
XFILLER_78_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14994_ _05891_ _05888_ net65 _05892_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__a211oi_2
X_16733_ a_l\[6\] net491 VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__nand2_1
XFILLER_81_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19521_ _10153_ _00571_ _00570_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__a21boi_2
X_13945_ _01888_ _04555_ _04846_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__o21a_1
XFILLER_35_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16664_ _07522_ _07532_ VGND VGND VPWR VPWR _07536_ sky130_fd_sc_hd__nand2_4
X_19452_ _10170_ _00637_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__nand2_1
X_13876_ _04780_ _04781_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__nand2_1
X_15615_ _06496_ _06433_ _06493_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__nand3_1
X_18403_ _09254_ _09256_ VGND VGND VPWR VPWR _09259_ sky130_fd_sc_hd__nand2_1
X_12827_ _03743_ _03750_ _03751_ VGND VGND VPWR VPWR _03756_ sky130_fd_sc_hd__nand3_2
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19383_ _10121_ net216 _10125_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__o21a_1
X_16595_ _07463_ _07464_ _07466_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__and3_1
X_18334_ _09176_ _09178_ _09180_ VGND VGND VPWR VPWR _09184_ sky130_fd_sc_hd__and3_1
XFILLER_50_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _09690_ _06426_ _06429_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__and3_1
XFILLER_91_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12758_ _03452_ _03531_ _03567_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__o22a_1
X_11709_ _02606_ _02641_ _02643_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__nand3_4
X_12689_ _03566_ net290 _03563_ _03615_ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__o211ai_4
X_18265_ net373 _09087_ net233 _09091_ VGND VGND VPWR VPWR _09111_ sky130_fd_sc_hd__o2bb2ai_1
X_15477_ _06345_ _06365_ _06367_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17216_ _08081_ _08078_ _08073_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__nand3_2
X_18196_ _09037_ _09038_ net458 _06401_ VGND VGND VPWR VPWR _09043_ sky130_fd_sc_hd__nand4_1
X_14428_ net723 net699 VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__nand2_1
Xmax_cap402 _02345_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_1
XFILLER_128_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17147_ _08012_ _08013_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__nand2_1
XFILLER_116_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14359_ _05102_ net142 _05261_ _05101_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__o211ai_4
Xmax_cap413 _09607_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_1
Xmax_cap468 _01754_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
X_17078_ _07830_ _07833_ _07944_ _07945_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__nand4_4
Xmax_cap457 _04260_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_12
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16029_ _06900_ _06902_ _06897_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__a21o_1
Xmax_cap479 net480 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__buf_6
XFILLER_69_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19719_ _00918_ _00922_ _00925_ _00921_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__o211a_1
XFILLER_53_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20425_ clknet_leaf_28_clk _00065_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20356_ net794 net53 VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__and2_1
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20287_ _01530_ _01531_ _01511_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__a21oi_1
X_11991_ _02861_ _02920_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__nand2_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10942_ net697 net691 net545 net538 VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__nand4_4
XFILLER_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13730_ _04633_ _04636_ _04631_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10873_ _09690_ net1183 VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__and2_1
X_13661_ _04566_ _04568_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__a21oi_4
X_15400_ _06247_ _06289_ _06248_ _06240_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__nand4_1
XFILLER_32_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16380_ _07240_ _07241_ _07247_ _07250_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__o2bb2ai_1
X_12612_ _03541_ net489 net665 _03539_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__nand4_1
X_13592_ _04488_ _04498_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_14_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12543_ _03469_ _03470_ _03465_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__a21o_1
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15331_ _06223_ _06224_ net719 net657 VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__nand4_4
XFILLER_24_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18050_ _08897_ net305 VGND VGND VPWR VPWR _08899_ sky130_fd_sc_hd__nor2_4
X_15262_ _06153_ _06155_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__nor2_1
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17001_ _07706_ _07708_ _07707_ VGND VGND VPWR VPWR _07871_ sky130_fd_sc_hd__o21a_1
X_12474_ _03394_ _03395_ net355 VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_78_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14213_ _05039_ _05081_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__nand2_1
X_11425_ _02361_ _02364_ _02356_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_78_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_7 _00352_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15193_ _06087_ _06088_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__nor2_1
XFILLER_125_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11356_ net967 net517 _02295_ _02296_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__a22oi_1
X_14144_ _05042_ _05045_ _05047_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_91_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18952_ _09773_ _09841_ _09842_ VGND VGND VPWR VPWR _09844_ sky130_fd_sc_hd__nand3_1
XFILLER_4_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ term_low\[21\] term_mid\[21\] _00687_ _00719_ VGND VGND VPWR VPWR _00762_
+ sky130_fd_sc_hd__o211ai_1
X_14075_ _04892_ _04898_ _04895_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__a21o_1
X_11287_ _02216_ _02219_ _02225_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__a21o_1
X_13026_ net136 _03605_ _03950_ _03951_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__nand4_4
X_17903_ _08734_ _08760_ VGND VGND VPWR VPWR _08762_ sky130_fd_sc_hd__xor2_1
X_18883_ _09639_ _09645_ _09642_ VGND VGND VPWR VPWR _09775_ sky130_fd_sc_hd__a21o_1
X_10238_ net794 net62 VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__and2_1
X_17834_ _09297_ _09679_ _08693_ VGND VGND VPWR VPWR _08695_ sky130_fd_sc_hd__o21ai_1
XFILLER_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17765_ _08614_ _08626_ _08627_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__a21oi_1
X_14977_ _05875_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__inv_2
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer19 net812 VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlymetal6s2s_1
X_16716_ _07580_ _07585_ _07583_ _07438_ VGND VGND VPWR VPWR _07587_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_89_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13928_ _04776_ _04808_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__nand2_1
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19504_ _00486_ _10160_ _00690_ _00684_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__o211ai_4
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17696_ _08552_ _08555_ _08556_ VGND VGND VPWR VPWR _08559_ sky130_fd_sc_hd__a21oi_1
X_16647_ _07514_ _07518_ _07517_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__o21ai_4
XFILLER_50_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13859_ _04763_ net318 _04761_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__nand3_2
X_19435_ _00614_ _00616_ _00610_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16578_ _07449_ _07448_ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__nand2_2
X_19366_ _09144_ _09384_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__nor2_1
XFILLER_22_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15529_ net628 net528 VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__nand2_1
X_18317_ _09163_ _09145_ VGND VGND VPWR VPWR _09165_ sky130_fd_sc_hd__nand2_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19297_ _10013_ _10016_ net898 VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_100_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18248_ _08898_ _09012_ _09003_ _09010_ VGND VGND VPWR VPWR _09095_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_30_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold502 p_hh\[25\] VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
X_18179_ net626 net754 VGND VGND VPWR VPWR _09026_ sky130_fd_sc_hd__nand2_1
XFILLER_143_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold524 term_high\[59\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _01655_ VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 term_high\[63\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap221 net223 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
X_20210_ _01351_ _01452_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__and2_1
XFILLER_143_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold579 term_high\[57\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 term_high\[52\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap254 _08753_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__clkbuf_1
Xmax_cap276 _09190_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_1
Xmax_cap265 net266 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
Xmax_cap287 _04626_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_4
X_20141_ _01366_ _01367_ _01374_ _01377_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__nand4_2
Xhold568 term_mid\[24\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
X_20072_ _01297_ _01301_ _01304_ _01299_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__o211a_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20408_ clknet_leaf_29_clk _00048_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfxtp_1
X_11210_ _02086_ _02090_ _02092_ _02074_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__a2bb2oi_1
X_12190_ _03036_ _03032_ _03035_ _03081_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__a22oi_4
XFILLER_135_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11141_ _02081_ _02083_ _09439_ _09592_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput66 net66 VGND VGND VPWR VPWR p[0] sky130_fd_sc_hd__buf_2
X_20339_ net793 net3 VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_73_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput88 net88 VGND VGND VPWR VPWR p[2] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR p[3] sky130_fd_sc_hd__buf_2
X_11072_ _02003_ _02009_ _02001_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__a21o_1
Xoutput77 net77 VGND VGND VPWR VPWR p[1] sky130_fd_sc_hd__buf_2
XFILLER_0_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15880_ net595 net531 VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__nand2_1
XFILLER_76_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14900_ net756 net750 net642 net640 VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__nand4_1
XFILLER_64_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14831_ _05712_ _05713_ _05726_ _05727_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__a22o_1
X_17550_ _08411_ _08412_ _08293_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_19_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ net561 net533 VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__nand2_1
X_11974_ _02890_ _02885_ _02889_ net323 _02907_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__o2111a_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14762_ _05661_ _05262_ _05260_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__nand3_4
X_10925_ _01870_ _01872_ _01868_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a21o_1
X_17481_ _08180_ _08183_ _08193_ _08345_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__o211ai_2
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13713_ _04604_ _04606_ _04611_ _04612_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__o2bb2ai_1
X_14693_ _05433_ net313 _05456_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__nand3_2
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16432_ _07301_ _07303_ _07172_ _07175_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__o2bb2ai_1
X_10856_ net793 net1223 VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__and2_1
X_13644_ _04549_ _04487_ _04548_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__nand3_4
X_19220_ _10069_ _10114_ net206 _10008_ VGND VGND VPWR VPWR _10118_ sky130_fd_sc_hd__o211ai_4
X_16363_ _09319_ _09581_ net1070 _07234_ _07233_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__o221ai_4
XFILLER_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19151_ net892 net562 net556 net776 VGND VGND VPWR VPWR _10043_ sky130_fd_sc_hd__a22oi_2
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10787_ _01782_ _01784_ _01810_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__o21bai_1
X_18102_ _08893_ _08946_ _08948_ VGND VGND VPWR VPWR _08951_ sky130_fd_sc_hd__nor3_1
X_13575_ _04389_ _04477_ _04483_ VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__a21oi_1
X_15314_ _06139_ _06205_ _06206_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__nand3b_2
X_16294_ _07165_ _07166_ net281 VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__and3_1
X_12526_ _03418_ _03457_ VGND VGND VPWR VPWR _03458_ sky130_fd_sc_hd__nand2_1
XFILLER_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19082_ _09904_ _09905_ _09966_ _09970_ VGND VGND VPWR VPWR _09973_ sky130_fd_sc_hd__nand4_2
X_18033_ _08865_ _08879_ _08881_ VGND VGND VPWR VPWR _08883_ sky130_fd_sc_hd__nand3_1
X_12457_ net665 net661 net499 net495 VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__nand4_2
X_15245_ _06137_ _06138_ _06080_ VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__nand3_1
X_11408_ net401 _02347_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__nand2_1
X_15176_ _06070_ _06072_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__nand2_1
XFILLER_99_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12388_ net460 _03319_ _03307_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__o211ai_4
X_14127_ _05004_ _05030_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nand2_1
X_11339_ _02277_ _02279_ _09460_ _09592_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_98_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19984_ net574 net568 net1043 net1098 VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__nand4_4
XFILLER_140_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14058_ _04962_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__nand2_2
X_18935_ _09824_ _09826_ VGND VGND VPWR VPWR _09827_ sky130_fd_sc_hd__nand2_1
XFILLER_67_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13009_ _03884_ _03885_ _03928_ _03930_ VGND VGND VPWR VPWR _03936_ sky130_fd_sc_hd__o2bb2ai_1
X_18866_ _04555_ _06605_ net619 net732 _09753_ VGND VGND VPWR VPWR _09758_ sky130_fd_sc_hd__o2111ai_4
XFILLER_95_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17817_ net555 net486 VGND VGND VPWR VPWR _08678_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18797_ _09210_ _09264_ _09684_ _09685_ VGND VGND VPWR VPWR _09689_ sky130_fd_sc_hd__o211ai_1
X_17748_ _08533_ _08535_ _08534_ VGND VGND VPWR VPWR _08611_ sky130_fd_sc_hd__a21bo_1
XFILLER_82_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17679_ _08541_ _08542_ VGND VGND VPWR VPWR _08543_ sky130_fd_sc_hd__and2_1
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20690_ clknet_3_4__leaf_clk _00330_ VGND VGND VPWR VPWR p_hl\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19418_ net588 net579 net835 net738 VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__nand4_1
X_19349_ _10092_ _10095_ _10098_ _10085_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_135_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold387 p_hh_pipe\[0\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 term_low\[6\] VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 p_ll\[7\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold398 mid_sum\[20\] VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
X_20124_ net731 net551 VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__nand2_1
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20055_ _01281_ _01282_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__nand2_1
XFILLER_86_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10710_ _01743_ _01744_ _01742_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__a21oi_1
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11690_ net658 net520 VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__nand2_1
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10641_ p_hl\[3\] p_lh\[3\] VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__nor2_1
XFILLER_10_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13360_ net772 net766 net701 net693 VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__nand4_2
X_10572_ net794 net1300 VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12311_ _03108_ _03104_ _03101_ _03105_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_127_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13291_ _04179_ _04202_ _04203_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__nand3b_1
X_12242_ net687 net483 net481 net692 VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__a22o_1
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15030_ net739 net733 net657 net651 VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__nand4_2
XFILLER_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12173_ _02789_ _02938_ _02939_ _03107_ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__a31o_1
X_16981_ _07695_ _07733_ _07846_ _07848_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__a2bb2oi_4
X_11124_ net686 net519 VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__nand2_1
X_15932_ _06789_ _06806_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__nor2_1
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11055_ _01955_ _01972_ net328 VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__a21oi_4
XFILLER_107_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18720_ net609 net743 net737 net619 VGND VGND VPWR VPWR _09605_ sky130_fd_sc_hd__a22oi_4
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15863_ _06582_ _06721_ _06713_ _06718_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18651_ _09445_ _09525_ _09524_ VGND VGND VPWR VPWR _09530_ sky130_fd_sc_hd__nand3_4
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15794_ _06596_ _06614_ _06615_ net382 VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__o2bb2ai_1
X_17602_ _08448_ _08453_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__nand2_1
X_18582_ net597 net759 net1001 net606 VGND VGND VPWR VPWR _09454_ sky130_fd_sc_hd__a22o_1
X_14814_ _05712_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__nand2_2
XFILLER_123_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11957_ _02737_ _02740_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__nand2_1
XFILLER_91_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ net565 net560 net500 net494 VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__and4_1
X_14745_ _05641_ _05551_ _05549_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__a21oi_1
X_10908_ net707 net947 net538 net713 VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a22o_1
X_17464_ _08316_ _08325_ _08327_ _08324_ VGND VGND VPWR VPWR _08330_ sky130_fd_sc_hd__o211a_1
X_16415_ _07284_ _07287_ _07154_ _07160_ _07288_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__o221ai_4
X_11888_ _02760_ net248 _02759_ _02796_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19203_ _10079_ _10081_ _10099_ VGND VGND VPWR VPWR _10100_ sky130_fd_sc_hd__o21ai_2
X_14676_ _05573_ _05575_ net745 net662 VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__nand4_4
X_17395_ _08254_ _08255_ _08240_ _08244_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__o211ai_1
X_10839_ net1373 net1341 _01854_ _01847_ net795 VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__o221a_1
X_13627_ _04511_ _04512_ _04530_ _04534_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_43_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16346_ _07212_ _07214_ _07215_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__nand3_1
X_13558_ net1133 _04463_ _04396_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__a21o_1
X_19134_ _10022_ _10012_ VGND VGND VPWR VPWR _10025_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16277_ net280 _07127_ _07143_ _07144_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__o2bb2ai_4
X_12509_ _03260_ b_h\[8\] net1019 VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__and3_1
X_19065_ _09926_ _09955_ VGND VGND VPWR VPWR _09956_ sky130_fd_sc_hd__nand2_1
X_18016_ net459 _06521_ _08837_ VGND VGND VPWR VPWR _08866_ sky130_fd_sc_hd__o21a_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13489_ _04345_ _04358_ _04353_ _04357_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__o2bb2ai_4
X_15228_ _06118_ _06119_ _06120_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__a21o_1
XFILLER_114_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15159_ _05996_ _06050_ _06051_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__and3_1
XFILLER_141_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19967_ _01143_ _01145_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__nand2_1
XFILLER_68_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18918_ _09656_ _09661_ _09659_ VGND VGND VPWR VPWR _09810_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_26_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19898_ _01017_ _01018_ _01022_ _01016_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__a22o_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18849_ _09688_ _09699_ VGND VGND VPWR VPWR _09741_ sky130_fd_sc_hd__nand2_1
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20742_ clknet_leaf_42_clk _00382_ VGND VGND VPWR VPWR p_ll\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20673_ clknet_leaf_5_clk _00313_ VGND VGND VPWR VPWR p_hl\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20107_ _01262_ _01277_ _01340_ _01341_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__a22oi_1
XFILLER_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20038_ _01086_ _01165_ _01175_ _01267_ _01266_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__o2111ai_4
X_12860_ _03710_ _03787_ _03788_ VGND VGND VPWR VPWR _03789_ sky130_fd_sc_hd__nand3_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11811_ _02728_ _02729_ _02745_ _02746_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__nand4_1
XFILLER_27_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _03717_ _03668_ _03662_ VGND VGND VPWR VPWR _03720_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_68_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _05301_ _05306_ _05303_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__a21bo_2
X_11742_ _02243_ net402 _02469_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11673_ net644 net546 net537 net1016 VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_81_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _05362_ _05363_ _05220_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16200_ _07071_ _07067_ _07065_ _07070_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__o211a_1
XFILLER_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17180_ _07812_ _07906_ _08045_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__a21o_2
X_13412_ _04321_ _04322_ _09177_ _09264_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_40_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ net794 net1262 VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__and2_1
X_14392_ _05290_ _05282_ VGND VGND VPWR VPWR _05295_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16131_ _06998_ _07001_ _06995_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__a21oi_1
X_13343_ _04211_ _04255_ net796 VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__a21oi_1
X_10555_ net793 net1221 VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__and2_1
X_10486_ _01645_ term_high\[49\] net796 VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__a21oi_1
X_16062_ _06936_ _06745_ _06934_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__and3_1
Xrebuffer292 _09171_ VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlymetal6s4s_1
X_13274_ _04181_ _04185_ a_h\[0\] net763 VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__and4_1
XFILLER_6_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer270 net1085 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
X_12225_ _03147_ _03153_ _03154_ VGND VGND VPWR VPWR _03159_ sky130_fd_sc_hd__nand3b_2
X_15013_ _05909_ _05910_ _05905_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__a21oi_1
X_12156_ _02829_ _02827_ _02828_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_9_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19821_ _01009_ _01011_ _01031_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__o21ai_2
X_11107_ _01996_ _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__nand2_1
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16964_ _07800_ _07801_ _07830_ _07831_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__o211a_2
X_12087_ _02999_ _03001_ _03013_ _03015_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__a22oi_4
X_19752_ _00861_ _00957_ _00958_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__nand3_2
X_15915_ net624 net505 VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__nand2_1
X_11038_ _01907_ _01911_ net466 VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__a21o_1
X_16895_ _07763_ _07746_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__nand2_1
XFILLER_77_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18703_ _09586_ _09580_ _09585_ VGND VGND VPWR VPWR _09587_ sky130_fd_sc_hd__a21oi_2
X_19683_ b_l\[8\] _00748_ net567 _00745_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__a31o_4
X_15846_ _06720_ _06721_ _06582_ VGND VGND VPWR VPWR _06725_ sky130_fd_sc_hd__a21o_1
XFILLER_92_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18634_ _09510_ _09474_ _09509_ VGND VGND VPWR VPWR _09511_ sky130_fd_sc_hd__and3_4
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15777_ _06587_ _06590_ net1051 VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__o21a_1
XFILLER_92_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18565_ _09432_ _09434_ _09435_ VGND VGND VPWR VPWR _09436_ sky130_fd_sc_hd__a21o_1
X_12989_ _03822_ _03827_ _03829_ net395 _03910_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__o2111ai_4
XFILLER_18_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17516_ _08209_ net416 _08290_ _08287_ _08378_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__a221o_1
X_18496_ net1124 net1146 net593 net585 VGND VGND VPWR VPWR _09360_ sky130_fd_sc_hd__nand4_1
X_14728_ _05628_ _05600_ _05627_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__nand3_2
X_17447_ _08311_ net448 _08303_ _08312_ VGND VGND VPWR VPWR _08313_ sky130_fd_sc_hd__o211ai_4
X_14659_ _05553_ _05557_ _05556_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17378_ _08094_ _08097_ net450 VGND VGND VPWR VPWR _08245_ sky130_fd_sc_hd__a21oi_1
X_19117_ _09976_ _09989_ VGND VGND VPWR VPWR _10007_ sky130_fd_sc_hd__nand2_2
XFILLER_9_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16329_ net629 net484 net480 a_l\[0\] VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__a22oi_1
X_19048_ net764 net575 VGND VGND VPWR VPWR _09939_ sky130_fd_sc_hd__nand2_1
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20725_ clknet_leaf_23_clk _00365_ VGND VGND VPWR VPWR p_lh\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20656_ clknet_leaf_12_clk _00296_ VGND VGND VPWR VPWR p_hh\[22\] sky130_fd_sc_hd__dfxtp_1
X_20587_ clknet_leaf_14_clk _00227_ VGND VGND VPWR VPWR p_hh_pipe\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10340_ term_low\[27\] term_mid\[27\] term_low\[26\] term_mid\[26\] VGND VGND VPWR
+ VPWR _01117_ sky130_fd_sc_hd__o211a_1
XFILLER_124_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10271_ _10083_ _10050_ net794 _10094_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__o211a_1
X_12010_ net247 _02942_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__o21ai_2
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone207 net1005 VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__clkbuf_16
Xclone218 net1017 VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__clkbuf_16
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13961_ _04856_ _04857_ _04860_ _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__a31o_1
X_16680_ _07507_ _07508_ _07546_ _07547_ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__a22o_1
X_15700_ _09231_ _09526_ _06536_ _06535_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__o31a_1
XFILLER_86_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12912_ _03814_ _03816_ _03836_ _03837_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__o211ai_4
XFILLER_47_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13892_ _04798_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__inv_2
XFILLER_0_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15631_ _06472_ _06490_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12843_ _03770_ _03735_ _03769_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__nand3_2
X_15562_ _06439_ _06442_ _06437_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__a21oi_1
X_12774_ _03702_ _03703_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__and2_1
X_18350_ _09112_ _09196_ _09197_ VGND VGND VPWR VPWR _09202_ sky130_fd_sc_hd__nand3_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11725_ _02657_ _02659_ _02648_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__nand3b_1
X_17301_ net584 net488 VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__nand2_2
X_18281_ _09113_ _09124_ _09125_ VGND VGND VPWR VPWR _09127_ sky130_fd_sc_hd__and3_1
X_15493_ _06359_ _06377_ _06379_ _06380_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__or4bb_1
X_14513_ _05318_ _05320_ _05298_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__o21ai_1
X_17232_ _09210_ _09668_ _08097_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__o21ai_2
X_14444_ net736 net677 VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__nand2_2
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11656_ _02587_ _02592_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__nand2_1
X_11587_ _02522_ net507 net1078 VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__nand3_1
X_17163_ _07893_ _07894_ _07896_ _07997_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__o2bb2a_1
X_10607_ net794 net1196 VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__and2_1
X_14375_ _05274_ _05275_ _05270_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10538_ net793 net1207 VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__and2_1
Xmax_cap617 net620 VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__buf_12
X_16114_ _06979_ _06987_ _06988_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__nand3_2
Xmax_cap606 net608 VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__buf_8
X_17094_ _07950_ _07956_ _07957_ VGND VGND VPWR VPWR _07963_ sky130_fd_sc_hd__nand3_4
X_13326_ net763 net710 _04236_ _04238_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a22o_1
XFILLER_10_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16045_ _06920_ _06914_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__nand2_2
Xmax_cap628 net629 VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_12
X_13257_ _04157_ _04158_ _04168_ _04170_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__or4bb_4
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap639 net640 VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__buf_12
X_10469_ term_mid\[47\] term_high\[47\] VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__xor2_1
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12208_ _03138_ _03139_ _03140_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_94_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13188_ _04104_ _04096_ _04103_ _04084_ _04082_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__o311a_1
X_12139_ _03068_ net268 _03071_ _02844_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__o2bb2ai_2
X_17996_ _08844_ _08845_ _08846_ VGND VGND VPWR VPWR _08847_ sky130_fd_sc_hd__o21ai_2
X_19804_ net735 net567 VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__nand2_1
X_16947_ _07644_ _07653_ _07810_ _07812_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__nand4_1
X_19735_ _00940_ _00942_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16878_ _07603_ _07606_ _07607_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__a21oi_2
XFILLER_65_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19666_ _00777_ _00823_ _00826_ _00778_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__a31oi_1
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15829_ _06700_ _06702_ _06689_ _06691_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__o211ai_1
X_18617_ _09485_ _09486_ VGND VGND VPWR VPWR _09492_ sky130_fd_sc_hd__nand2_1
XFILLER_53_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19597_ _00596_ _00597_ _00595_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__a21oi_1
X_18548_ _09414_ _09415_ VGND VGND VPWR VPWR _09418_ sky130_fd_sc_hd__nand2_1
XFILLER_18_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20510_ clknet_leaf_32_clk _00150_ VGND VGND VPWR VPWR term_low\[5\] sky130_fd_sc_hd__dfxtp_1
X_18479_ _09338_ _09327_ VGND VGND VPWR VPWR _09342_ sky130_fd_sc_hd__nand2_1
X_20441_ clknet_leaf_28_clk _00081_ VGND VGND VPWR VPWR term_high\[33\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20372_ clknet_leaf_52_clk _00012_ VGND VGND VPWR VPWR b_l\[12\] sky130_fd_sc_hd__dfxtp_4
XFILLER_134_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11510_ _02342_ _02341_ _02340_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__o21ai_1
X_12490_ _03151_ _03420_ VGND VGND VPWR VPWR _03422_ sky130_fd_sc_hd__or2_1
X_20708_ clknet_leaf_41_clk net135 VGND VGND VPWR VPWR p_lh\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20639_ clknet_leaf_26_clk _00279_ VGND VGND VPWR VPWR p_hh\[5\] sky130_fd_sc_hd__dfxtp_1
Xwire136 _03607_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_6
X_11441_ _02376_ _02377_ net681 net517 VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__nand4_2
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11372_ _02268_ _02269_ _02309_ _02310_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__nand4_2
XFILLER_50_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14160_ _05059_ _05060_ _05051_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__and3_1
XFILLER_124_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13111_ _03953_ _04035_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__nand2_1
X_10323_ _00913_ _00924_ net794 VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__o21ai_1
X_14091_ _04986_ _04989_ _04982_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__a21o_1
XFILLER_140_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10254_ _09690_ net1312 VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13042_ _03903_ _03964_ _03967_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__a21oi_2
X_17850_ _08708_ _08710_ VGND VGND VPWR VPWR _08711_ sky130_fd_sc_hd__nand2_1
X_10185_ net897 VGND VGND VPWR VPWR _09199_ sky130_fd_sc_hd__inv_12
XFILLER_59_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16801_ net584 net572 net513 net506 VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__nand4_2
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17781_ _08641_ _08642_ VGND VGND VPWR VPWR _08643_ sky130_fd_sc_hd__nand2_1
X_19520_ _10152_ _10153_ _00570_ _00571_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__nand4_4
X_14993_ _05890_ _05883_ _05881_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__and3_1
X_16732_ net608 net488 VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__nand2_1
XFILLER_75_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13944_ _04844_ _04845_ _04846_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__a21oi_1
X_16663_ _07524_ _07527_ net970 VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__nand3_2
X_19451_ b_l\[3\] net548 VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__nand2_1
X_13875_ net734 net703 net699 net741 VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__a22oi_2
XFILLER_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15614_ _06462_ _06494_ _06495_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__nand3_2
X_18402_ _09231_ _09242_ net805 _09248_ _09250_ VGND VGND VPWR VPWR _09258_ sky130_fd_sc_hd__o311a_1
X_12826_ _03754_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__inv_2
X_19382_ _10121_ net216 _10125_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16594_ _07324_ _07327_ _07326_ VGND VGND VPWR VPWR _07466_ sky130_fd_sc_hd__a21boi_1
X_18333_ _09172_ _09131_ _09083_ _09179_ VGND VGND VPWR VPWR _09183_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_17_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _06425_ _06428_ _06410_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__a21o_1
X_12757_ _03532_ _03569_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__nand2_1
XFILLER_147_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11708_ _02639_ _02640_ _02605_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__a21oi_1
X_12688_ _03615_ _03617_ _03565_ VGND VGND VPWR VPWR _03618_ sky130_fd_sc_hd__nand3b_2
X_18264_ _09090_ _09024_ _09088_ net373 VGND VGND VPWR VPWR _09110_ sky130_fd_sc_hd__a31o_1
X_15476_ _06365_ _06345_ net795 VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__o21ai_1
X_11639_ _02456_ _02451_ _02455_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_96_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17215_ _07916_ _08080_ _08079_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__a21oi_2
X_18195_ _08955_ net336 VGND VGND VPWR VPWR _09042_ sky130_fd_sc_hd__or2_1
X_14427_ net727 net695 VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__nand2_1
X_17146_ _08009_ _08011_ _08014_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_96_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _05100_ _05256_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__and2_4
XFILLER_128_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire692 net696 VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__buf_12
X_13309_ net787 net933 VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__nand2_1
Xmax_cap425 _05576_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_2
X_17077_ _07936_ _07942_ _07940_ VGND VGND VPWR VPWR _07946_ sky130_fd_sc_hd__o21ai_1
Xmax_cap447 _09605_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_4
X_14289_ net724 net703 net699 net727 VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__a22o_2
Xmax_cap458 _04259_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__buf_6
X_16028_ _09144_ _09613_ _06794_ _06901_ _06900_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__o221ai_2
XFILLER_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17979_ net338 net306 _08830_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__o21a_1
XFILLER_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19718_ _00801_ _00802_ _00799_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__a21oi_2
X_19649_ _00702_ _00850_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20424_ clknet_leaf_28_clk _00064_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20355_ net794 net52 VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__and2_1
XFILLER_122_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20286_ _09362_ _09373_ _01529_ _01531_ _01511_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__o311a_1
XFILLER_121_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11990_ _02925_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__inv_2
X_10941_ net700 net693 VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__nand2_8
XFILLER_17_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13660_ _04461_ _04395_ _04462_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__a21o_4
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10872_ _09690_ net1155 VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__and2_1
X_12611_ _03539_ _03541_ _09471_ _09646_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13591_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12542_ _03469_ _03470_ _03465_ VGND VGND VPWR VPWR _03474_ sky130_fd_sc_hd__a21oi_1
X_15330_ net726 net722 net871 net643 VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__nand4_2
X_12473_ _03401_ _03403_ _03402_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a21o_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15261_ _06150_ _06152_ net719 net1019 VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__nand4_1
X_17000_ _07706_ _07708_ _07707_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__o21ai_2
X_11424_ net658 net652 net546 net539 VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_78_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14212_ _05114_ _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__nand2_2
XANTENNA_8 _00424_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15192_ _06086_ _06083_ _06085_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__and3_1
X_11355_ _02159_ _02293_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__nand2_1
X_14143_ _05042_ _05046_ _05047_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__nand3b_1
X_11286_ _02222_ _02223_ _02216_ _02219_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_91_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18951_ _09773_ _09842_ VGND VGND VPWR VPWR _09843_ sky130_fd_sc_hd__nand2_1
X_14074_ _04974_ _04977_ _04978_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__o21ai_2
X_10306_ _00709_ _00730_ _00741_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__o21a_1
XFILLER_140_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13025_ _03602_ _03704_ _03790_ _03875_ VGND VGND VPWR VPWR _03952_ sky130_fd_sc_hd__nand4b_4
X_17902_ _09319_ _09679_ _08728_ _08733_ _08760_ VGND VGND VPWR VPWR _08761_ sky130_fd_sc_hd__o311a_1
X_10237_ net794 net61 VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__and2_1
XFILLER_121_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18882_ _09640_ _09641_ _09639_ VGND VGND VPWR VPWR _09774_ sky130_fd_sc_hd__a21oi_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17833_ net900 net473 _08691_ _08693_ VGND VGND VPWR VPWR _08694_ sky130_fd_sc_hd__a22o_1
X_17764_ _08614_ _08626_ net795 VGND VGND VPWR VPWR _08627_ sky130_fd_sc_hd__o21ai_1
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14976_ _09384_ _09417_ _05756_ _05754_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__o31a_1
X_16715_ _07580_ _07585_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__nand2_4
X_13927_ _04777_ _04795_ _04796_ _04800_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__a31o_1
X_19503_ _00684_ _00686_ _00689_ _00489_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_89_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17695_ _08481_ _08553_ net1093 net478 _08552_ VGND VGND VPWR VPWR _08558_ sky130_fd_sc_hd__o2111ai_2
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19434_ _00616_ net718 net887 _00614_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__and4_1
X_16646_ _06999_ _07513_ _07512_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__o21ai_2
XFILLER_90_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13858_ _04763_ net318 _04761_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__and3_1
XFILLER_23_808 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16577_ _09166_ _09679_ _07444_ _07445_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__o211ai_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ net659 net486 b_h\[13\] net920 VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__a22o_1
X_13789_ _04475_ _04574_ _04575_ _04692_ _04694_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__a41o_1
X_19365_ _10071_ _00538_ _00539_ _00540_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_33_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ net623 net540 VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__nand2_1
X_18316_ _09140_ _09141_ _09162_ VGND VGND VPWR VPWR _09164_ sky130_fd_sc_hd__o21ai_4
X_19296_ _00462_ _00464_ _00453_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_100_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18247_ _09091_ net233 net373 _09087_ VGND VGND VPWR VPWR _09094_ sky130_fd_sc_hd__o211ai_2
XFILLER_135_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15459_ _06315_ _06314_ _06349_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__a21oi_1
Xmax_cap200 _02321_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__buf_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18178_ net630 net749 VGND VGND VPWR VPWR _09025_ sky130_fd_sc_hd__nand2_1
Xmax_cap211 _04685_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__buf_1
XFILLER_144_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold514 _01672_ VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 p_hh\[1\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ _07896_ _07997_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__nor2_1
Xhold536 p_hh\[31\] VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap233 _09089_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__buf_1
Xhold503 mid_sum\[11\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap222 _06355_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
Xhold558 term_high\[61\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold569 p_lh\[30\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap277 _09044_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__buf_4
Xmax_cap266 _04074_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
Xhold547 p_ll\[31\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ _01366_ _01367_ _01374_ _01377_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__a22o_1
XFILLER_103_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap299 _09697_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_1
Xmax_cap288 _04564_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
XFILLER_106_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20071_ _01217_ _01222_ _01219_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o21ai_2
XFILLER_100_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20407_ clknet_leaf_47_clk _00047_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11140_ net678 net671 net547 net538 VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__nand4_2
XFILLER_107_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20338_ net793 net2 VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__and2_1
XFILLER_122_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput67 net67 VGND VGND VPWR VPWR p[10] sky130_fd_sc_hd__buf_2
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11071_ _02014_ _02001_ _02013_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__nand3_2
Xoutput89 net89 VGND VGND VPWR VPWR p[30] sky130_fd_sc_hd__buf_2
X_20269_ _01472_ _01469_ _01473_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__a21boi_1
Xoutput78 net78 VGND VGND VPWR VPWR p[20] sky130_fd_sc_hd__buf_2
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14830_ _05714_ _05726_ _05727_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__nand3_2
XFILLER_56_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ net570 net529 VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__nand2_1
X_11973_ _02890_ _02885_ _02889_ _02907_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__o211ai_1
X_14761_ _05407_ _05408_ _05532_ _05533_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__nand4_4
X_10924_ net702 net697 net545 net538 VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__nand4_2
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17480_ _08192_ _08344_ _08343_ VGND VGND VPWR VPWR _08346_ sky130_fd_sc_hd__o21bai_1
X_13712_ _04604_ _04606_ _04617_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__nand3_1
X_14692_ _05589_ _05590_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__nand2_1
X_10855_ net793 net1278 VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__and2_1
X_16431_ _07171_ _07301_ _07174_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__nand3_1
XFILLER_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13643_ _04548_ _04487_ _04549_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__and3_4
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16362_ _07233_ _07235_ _07229_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__a21o_1
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13574_ _04314_ _04476_ _04388_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__a21oi_1
X_19150_ net776 net556 VGND VGND VPWR VPWR _10042_ sky130_fd_sc_hd__nand2_1
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10786_ net442 _01789_ _01794_ _01803_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__nand4_1
X_18101_ _08946_ _08948_ VGND VGND VPWR VPWR _08950_ sky130_fd_sc_hd__or2_1
X_12525_ net292 _03453_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__o21ai_2
XFILLER_9_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15313_ _06205_ _06206_ _06139_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__a21bo_1
X_16293_ _07166_ _07165_ _07033_ _07034_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__o2bb2ai_4
X_19081_ _09906_ _09971_ VGND VGND VPWR VPWR _09972_ sky130_fd_sc_hd__nand2_1
XFILLER_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12456_ net665 net661 net495 VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__nand3_1
X_18032_ _08879_ _08881_ _08865_ VGND VGND VPWR VPWR _08882_ sky130_fd_sc_hd__a21o_1
X_15244_ _06137_ _06138_ _06080_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__a21o_1
X_11407_ _02243_ _02345_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__nand2_2
X_12387_ _03313_ _03315_ _03309_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__a21o_1
X_15175_ _06066_ _06067_ _06068_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__nand3_2
XFILLER_141_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11338_ net664 net658 net547 net539 VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__nand4_1
X_14126_ _05030_ _05006_ _05004_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__nand3b_1
XFILLER_141_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19983_ net574 net568 net1043 net1095 VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__and4_1
X_11269_ net464 _02201_ net361 _02199_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__o211ai_1
X_14057_ _04959_ _04961_ _04822_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__nand3_1
X_18934_ _09819_ _09814_ _09810_ _09818_ VGND VGND VPWR VPWR _09826_ sky130_fd_sc_hd__o211ai_4
X_13008_ _03884_ _03885_ _03929_ _03931_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__nand4_1
X_18865_ _04555_ _06605_ net619 net732 _09753_ VGND VGND VPWR VPWR _09757_ sky130_fd_sc_hd__o2111a_4
XFILLER_94_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17816_ net960 net999 VGND VGND VPWR VPWR _08677_ sky130_fd_sc_hd__nand2_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18796_ _09687_ _09678_ _09686_ VGND VGND VPWR VPWR _09688_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_38_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17747_ _08471_ _08473_ _08607_ _08608_ VGND VGND VPWR VPWR _08610_ sky130_fd_sc_hd__nand4_1
X_14959_ _05850_ _05853_ _05855_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__nand3_1
XFILLER_35_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17678_ _08538_ _08466_ _08537_ VGND VGND VPWR VPWR _08542_ sky130_fd_sc_hd__nand3_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16629_ net950 net502 _07497_ _07499_ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19417_ _04555_ _06985_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__nor2_1
XFILLER_62_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19348_ _10085_ _10098_ _10095_ _10092_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__o2bb2a_1
XPHY_EDGE_ROW_99_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19279_ _10179_ _10162_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__nand2_4
XFILLER_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold366 p_ll_pipe\[3\] VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 p_ll\[24\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold388 p_ll\[5\] VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold399 p_ll_pipe\[13\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20123_ _01293_ _01297_ _01295_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__o21ai_1
XFILLER_133_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20054_ net568 net1013 net1044 net1097 VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__nand4_1
XFILLER_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ _01685_ _01684_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__and2b_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10571_ net794 net1283 VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__and2_1
X_12310_ _03239_ _03238_ _03240_ VGND VGND VPWR VPWR _03244_ sky130_fd_sc_hd__and3_4
X_13290_ _04202_ _04203_ _04180_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__a21o_1
XFILLER_6_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12241_ net687 net481 VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__nand2_1
XFILLER_107_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12172_ _09177_ _09679_ _02941_ VGND VGND VPWR VPWR _03107_ sky130_fd_sc_hd__nor3_1
X_11123_ net967 net525 net519 net691 VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__a22o_1
X_16980_ _07735_ _07846_ _07848_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__nand3_2
X_15931_ _06660_ _06788_ _06806_ _06807_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__o211a_1
X_11054_ _01968_ _01956_ _01967_ _01951_ _01950_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__a32oi_1
XFILLER_110_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18650_ _09511_ _09521_ _09446_ _09523_ VGND VGND VPWR VPWR _09529_ sky130_fd_sc_hd__o211ai_4
X_15862_ _06538_ _06578_ _06579_ _06580_ _06721_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__o41a_1
X_17601_ _08353_ _08446_ _08447_ _08373_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__a31oi_1
XFILLER_67_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15793_ _06670_ _06671_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__nand2_1
XFILLER_92_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18581_ net597 net759 VGND VGND VPWR VPWR _09453_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14813_ net720 net690 _05710_ _05711_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__a22o_1
XFILLER_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11956_ _02733_ _02736_ _02739_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__o21ai_2
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17532_ _08309_ _08395_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__nand2_1
X_14744_ _05463_ _05550_ _05639_ _05640_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__a22o_1
XFILLER_17_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10907_ net544 net540 VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__nand2_8
X_17463_ _08324_ _08326_ _08327_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__a21o_1
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16414_ _07218_ _07220_ _07285_ _07286_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__a22o_1
X_11887_ _02759_ _02796_ _02760_ net248 VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__o2bb2ai_1
X_19202_ _10092_ _10095_ _10098_ VGND VGND VPWR VPWR _10099_ sky130_fd_sc_hd__o21ai_2
X_14675_ _09264_ _09482_ _05572_ _05574_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__o22ai_2
X_17394_ _08240_ _08244_ _08254_ _08255_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__o2bb2ai_1
X_10838_ p_hl\[30\] p_lh\[30\] p_hl\[31\] net1377 VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__a22o_1
XFILLER_60_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13626_ _04530_ _04534_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16345_ _07206_ _07211_ _07207_ _07216_ VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__a31oi_1
X_10769_ p_hl\[20\] p_lh\[20\] p_hl\[21\] p_lh\[21\] VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__a22o_1
X_13557_ _04463_ _04395_ net1133 VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__nand3_1
X_19133_ _09253_ _09264_ _10017_ _10019_ VGND VGND VPWR VPWR _10024_ sky130_fd_sc_hd__o211ai_2
X_16276_ _07127_ net280 _07146_ _07148_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_117_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12508_ _03435_ _03436_ _03427_ VGND VGND VPWR VPWR _03440_ sky130_fd_sc_hd__nand3_4
X_13488_ _04366_ _04333_ _04364_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__a21oi_4
X_19064_ _09937_ _09938_ _09944_ _09945_ VGND VGND VPWR VPWR _09955_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12439_ _03369_ _03370_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__nand2_1
X_18015_ _08863_ _08864_ VGND VGND VPWR VPWR _08865_ sky130_fd_sc_hd__nand2_4
X_15227_ _06118_ _06119_ _06121_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__nand3_4
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15158_ _05998_ _06048_ _05997_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__a21o_1
X_19966_ _01127_ _01131_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__nor2_1
X_14109_ net758 net752 net676 net670 VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__nand4_4
X_15089_ _05986_ _05985_ net65 VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__a21oi_1
X_18917_ _09656_ _09661_ _09659_ VGND VGND VPWR VPWR _09809_ sky130_fd_sc_hd__a21o_1
X_19897_ net742 net735 net1013 net556 _01109_ VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__a41o_1
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18848_ _09619_ _09598_ net335 VGND VGND VPWR VPWR _09740_ sky130_fd_sc_hd__a21boi_1
XFILLER_103_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18779_ _09667_ _09669_ VGND VGND VPWR VPWR _09670_ sky130_fd_sc_hd__nand2_1
X_20741_ clknet_leaf_41_clk _00381_ VGND VGND VPWR VPWR p_ll\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_733 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20672_ clknet_leaf_40_clk _00312_ VGND VGND VPWR VPWR p_hl\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_21_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_70_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20106_ _09253_ _01194_ _09384_ _01193_ _01339_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__o311ai_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20037_ _01262_ _01263_ net203 VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__a21o_1
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11810_ _02745_ _02746_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__nand2_1
X_12790_ _03661_ _03667_ _03717_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__o21ai_2
XFILLER_27_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _02573_ _02675_ _02676_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__nand3_1
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11672_ net644 net546 VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__nand2_1
X_14460_ _05138_ _05356_ _05357_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_81_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13411_ net751 net1076 net705 net757 VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a22o_4
XTAP_TAPCELL_ROW_40_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ net794 net1276 VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__and2_1
X_14391_ _05280_ _05281_ _05288_ _05289_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_40_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10554_ net793 net1281 VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__and2_1
X_16130_ _06996_ _06997_ _07004_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__a21o_1
X_13342_ _04253_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__nand2_1
XFILLER_10_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10485_ _01641_ _01642_ _01636_ _01635_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__a31o_1
X_16061_ _06743_ _06744_ _06934_ _06936_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__o211ai_2
X_13273_ _01860_ net805 net763 _04181_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__o211ai_1
Xrebuffer271 _04472_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__buf_2
Xrebuffer260 b_l\[0\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd1_1
X_12224_ _03157_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__inv_2
XFILLER_5_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15012_ _05908_ net642 net745 _05907_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__nand4_4
X_12155_ net177 _03089_ _03088_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__o21ai_2
XFILLER_123_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19820_ _01012_ _01028_ _01030_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__nand3_1
X_11106_ _02034_ _02035_ net363 VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__nand3_1
X_19751_ _00865_ _00866_ _00953_ _00955_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__a22o_1
X_16963_ _07800_ _07801_ _07831_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__o21ai_2
X_12086_ _03005_ _03018_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__nand2_1
XFILLER_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18702_ _09443_ _09576_ _09577_ _09437_ VGND VGND VPWR VPWR _09586_ sky130_fd_sc_hd__a31oi_2
X_11037_ net712 net1018 VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__nand2_1
X_15914_ net628 net502 VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__nand2_1
X_16894_ _07742_ _07744_ _07760_ _07762_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__o211ai_1
X_19682_ _00878_ _00880_ _00734_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__nand3_2
X_15845_ _06713_ _06718_ _06721_ _06582_ VGND VGND VPWR VPWR _06724_ sky130_fd_sc_hd__o211ai_1
XFILLER_77_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18633_ net301 _09496_ _09506_ _09507_ VGND VGND VPWR VPWR _09510_ sky130_fd_sc_hd__o2bb2ai_1
X_18564_ _09303_ _09299_ _09191_ _09306_ VGND VGND VPWR VPWR _09435_ sky130_fd_sc_hd__a22oi_4
X_15776_ _06587_ _06590_ net1051 VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__o21ai_2
X_17515_ _08209_ net416 _08290_ _08287_ _08378_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__a221oi_2
X_12988_ _03827_ _03911_ _03910_ net395 VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__o211a_1
X_11939_ net679 net1048 net511 net508 net438 VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__a41o_1
X_18495_ net1123 net1146 net593 net585 VGND VGND VPWR VPWR _09359_ sky130_fd_sc_hd__and4_1
X_14727_ _05606_ _05607_ _05622_ _05625_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__a22o_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17446_ _08308_ _08310_ _09286_ _09646_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__o2bb2ai_2
X_14658_ _05553_ _05554_ net761 net642 VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__o211a_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17377_ _08198_ _08242_ _08241_ _08239_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__o211ai_2
X_13609_ net777 net673 VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__nand2_1
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16328_ _07193_ _07201_ _07188_ _07200_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__o211ai_4
Xclkbuf_leaf_12_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_99_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19116_ _09870_ _09974_ _09975_ _09977_ _09987_ VGND VGND VPWR VPWR _10006_ sky130_fd_sc_hd__a32oi_4
XFILLER_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14589_ _05471_ _05473_ _05486_ _05487_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__o211ai_1
XFILLER_146_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16259_ _07129_ net505 net607 VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__nand3_1
X_19047_ net410 _09935_ _09936_ VGND VGND VPWR VPWR _09938_ sky130_fd_sc_hd__nand3_4
XFILLER_141_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19949_ _01160_ _01162_ _01086_ _01171_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__a31oi_1
XFILLER_101_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20724_ clknet_3_4__leaf_clk _00364_ VGND VGND VPWR VPWR p_lh\[26\] sky130_fd_sc_hd__dfxtp_1
X_20655_ clknet_leaf_11_clk _00295_ VGND VGND VPWR VPWR p_hh\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire318 _04728_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_2
XFILLER_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20586_ clknet_leaf_14_clk _00226_ VGND VGND VPWR VPWR p_hh_pipe\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10270_ _10050_ _10072_ term_low\[16\] net1316 VGND VGND VPWR VPWR _10094_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone219 net647 VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13960_ _04791_ _04792_ _04788_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a21boi_1
XFILLER_86_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12911_ _03838_ _03818_ VGND VGND VPWR VPWR _03839_ sky130_fd_sc_hd__nand2_2
X_15630_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__inv_2
XFILLER_74_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13891_ _04795_ _04796_ _04777_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__nand3_2
XFILLER_104_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12842_ _03769_ _03770_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__nand2_1
X_15561_ net1070 _06441_ net1120 net540 _06439_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__o2111ai_2
X_12773_ _03700_ _03701_ _03610_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__nand3_1
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11724_ _02657_ _02658_ _02648_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__o21bai_1
X_17300_ _08108_ _08110_ VGND VGND VPWR VPWR _08167_ sky130_fd_sc_hd__nand2_1
XFILLER_70_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18280_ _09124_ _09125_ _09113_ VGND VGND VPWR VPWR _09126_ sky130_fd_sc_hd__a21oi_2
XFILLER_42_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15492_ _06378_ _06379_ _06381_ _06359_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14512_ _05324_ _05180_ _05371_ _05328_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__o22ai_2
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11655_ net712 net983 net463 _02591_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a31o_1
X_17231_ _09210_ _09668_ _08097_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__o21a_1
X_14443_ _05207_ _05344_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__nand2_1
XFILLER_80_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17162_ net795 _08029_ _08030_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__and3_1
X_11586_ net1078 net681 net510 net507 VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__nand4_4
X_10606_ net794 net1230 VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__and2_1
X_14374_ _09220_ _09493_ _02613_ net805 _05274_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__o221ai_2
X_10537_ net793 net1240 VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__and2_1
X_16113_ _06979_ _06987_ _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__and3_1
X_17093_ _07749_ _07752_ _07958_ _07960_ _07755_ VGND VGND VPWR VPWR _07962_ sky130_fd_sc_hd__o221a_1
X_13325_ _04183_ _04235_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__nand2_1
Xmax_cap618 net619 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_12_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10468_ net796 _01629_ net140 VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__nor3_1
X_16044_ _06911_ _06912_ _06916_ _06894_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__a22o_1
Xmax_cap629 a_l\[1\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_8
X_13256_ _04157_ _04158_ _04168_ _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_110_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12207_ _03140_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10399_ _01570_ _01565_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__nand2_1
X_13187_ _04082_ _04084_ _04105_ _04106_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__a22o_1
X_12138_ net399 _02844_ _03070_ _02843_ VGND VGND VPWR VPWR _03073_ sky130_fd_sc_hd__o211a_1
XFILLER_97_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17995_ _08843_ _08835_ _08842_ VGND VGND VPWR VPWR _08846_ sky130_fd_sc_hd__nand3_1
X_19803_ net574 net731 VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__nand2_1
XFILLER_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16946_ _07644_ _07810_ _07812_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__nand3_2
X_12069_ net357 VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_19734_ _00793_ _00811_ _00809_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__a21o_1
X_19665_ _00865_ _00866_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_125_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16877_ _07603_ _07606_ _07607_ VGND VGND VPWR VPWR _07747_ sky130_fd_sc_hd__a21o_1
XFILLER_65_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18616_ _09155_ _09286_ _09371_ _09481_ _09480_ VGND VGND VPWR VPWR _09491_ sky130_fd_sc_hd__o221ai_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15828_ _06689_ _06691_ _06698_ _06699_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__o2bb2ai_1
X_19596_ _00790_ _00792_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__nor2_2
X_15759_ _06637_ _06508_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__nand2_1
X_18547_ _09414_ _09415_ VGND VGND VPWR VPWR _09416_ sky130_fd_sc_hd__nor2_1
X_18478_ _09334_ _09335_ _09330_ VGND VGND VPWR VPWR _09341_ sky130_fd_sc_hd__a21o_1
X_17429_ _08292_ _08294_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__nand2_2
X_20440_ clknet_leaf_29_clk _00080_ VGND VGND VPWR VPWR term_high\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20371_ clknet_leaf_52_clk _00011_ VGND VGND VPWR VPWR b_l\[11\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_31_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload50 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinv_8
XFILLER_115_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20707_ clknet_leaf_35_clk _00347_ VGND VGND VPWR VPWR p_lh\[9\] sky130_fd_sc_hd__dfxtp_2
X_20638_ clknet_leaf_26_clk _00278_ VGND VGND VPWR VPWR p_hh\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11440_ _02376_ _02377_ net681 net517 VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__and4_1
Xwire137 _08620_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
X_11371_ _02266_ _02267_ _02309_ _02310_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__a22o_1
Xwire159 _08007_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
X_20569_ clknet_leaf_7_clk _00209_ VGND VGND VPWR VPWR mid_sum\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13110_ _03950_ _03952_ _03951_ _04034_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__a31oi_2
X_14090_ _09155_ _09504_ _04893_ _04988_ _04986_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__o221ai_2
X_10322_ term_low\[24\] net1365 _00859_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__a21o_1
X_13041_ net634 net825 net885 net641 VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__a22oi_4
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10253_ _09690_ net1173 VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10184_ net1045 VGND VGND VPWR VPWR _09188_ sky130_fd_sc_hd__clkinv_8
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16800_ net578 net506 VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__nand2_2
X_17780_ _08632_ _08633_ _08638_ _08640_ VGND VGND VPWR VPWR _08642_ sky130_fd_sc_hd__nand4_2
X_16731_ _09210_ _09646_ VGND VGND VPWR VPWR _07602_ sky130_fd_sc_hd__nor2_1
XFILLER_93_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14992_ _05889_ _05884_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__and2_1
X_13943_ _04847_ _04848_ _04840_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__nand3_1
X_16662_ _07524_ _07528_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__nand2_1
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19450_ net765 net556 VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__nand2_1
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13874_ net741 net701 VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__nand2_1
X_16593_ _07327_ _07324_ _09624_ _07325_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__o2bb2ai_1
X_15613_ _06489_ _06490_ _06472_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__a21o_1
X_18401_ _09250_ _09251_ _09248_ VGND VGND VPWR VPWR _09257_ sky130_fd_sc_hd__a21oi_1
X_12825_ _03753_ _03742_ _03752_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__nand3_2
X_19381_ _00560_ _10159_ _00559_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__nand3_2
X_15544_ _06423_ _06424_ _06406_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__a21o_1
X_18332_ _09173_ _09174_ net232 VGND VGND VPWR VPWR _09182_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_120_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _03681_ _03684_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__o21ai_1
XFILLER_42_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11707_ _02606_ _02643_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__nand2_1
X_18263_ net797 _09108_ _09109_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__nor3_1
X_12687_ _03563_ _03566_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__nand2_1
X_15475_ _06341_ _06343_ _06365_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__a21oi_1
XFILLER_147_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11638_ _02451_ _02456_ _01871_ _02338_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_96_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _07936_ _07941_ _07916_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__o21a_1
X_18194_ _08955_ net336 VGND VGND VPWR VPWR _09041_ sky130_fd_sc_hd__nor2_1
X_14426_ _05327_ _05179_ _05326_ net1056 VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__nand4_4
X_17145_ _07857_ net472 a_l\[2\] _07855_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_96_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14357_ _05098_ _05255_ _05256_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__o21ai_2
Xmax_cap404 _01924_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_2
X_11569_ _02501_ _02503_ _09482_ _09592_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__o2bb2ai_1
X_13308_ net784 net933 VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__nand2_1
Xwire693 net696 VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__buf_6
Xmax_cap426 _05567_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_4
X_17076_ _07918_ _07937_ _07939_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__nand3_1
Xmax_cap448 _08307_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_2
Xmax_cap459 _04134_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__buf_12
X_14288_ net727 net724 net703 net699 VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__nand4_1
X_16027_ _06794_ _06901_ net624 net502 _06900_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__o2111ai_4
XFILLER_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13239_ net713 net710 _04133_ _04141_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__a41o_1
XFILLER_41_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_71_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17978_ net338 net306 net797 VGND VGND VPWR VPWR _08830_ sky130_fd_sc_hd__a21oi_1
X_16929_ _07667_ _07672_ _07669_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__a21oi_1
X_19717_ _00801_ _00802_ _00799_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__a21o_1
XFILLER_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19648_ _00549_ _00703_ _00701_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__o21ai_2
XFILLER_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19579_ _00643_ _00667_ _00669_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__nand3_1
XFILLER_37_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_80_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20423_ clknet_leaf_28_clk _00063_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20354_ net794 net51 VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__and2_1
XFILLER_88_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20285_ b_l\[14\] net548 net716 net551 VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__a22o_1
XFILLER_96_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10940_ net691 net947 VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__nand2_2
XFILLER_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10871_ net793 net1333 VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_119_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12610_ _03537_ _03538_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__nand2_2
X_13590_ _04492_ _04495_ _04497_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_14_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12541_ _03471_ _03470_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__nand2_1
XFILLER_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12472_ _03401_ _03403_ _03402_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__a21oi_1
X_15260_ _06150_ _06152_ net719 net1019 VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__and4_1
X_11423_ net658 net652 net539 VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__nand3_2
X_14211_ _05109_ _05112_ net714 b_l\[15\] VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__nand4_1
XANTENNA_9 _00434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15191_ _06085_ _06086_ _06083_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_128_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11354_ net681 net1061 net525 net519 VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__nand4_2
X_14142_ net714 net721 VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__nand2_1
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11285_ _02216_ _02219_ _02222_ _02223_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_91_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18950_ _09791_ _09792_ _09835_ _09837_ VGND VGND VPWR VPWR _09842_ sky130_fd_sc_hd__a22o_1
X_14073_ _04974_ _04975_ _04973_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__o21bai_4
X_10305_ _00709_ _00730_ net797 VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17901_ _08758_ _08759_ VGND VGND VPWR VPWR _08760_ sky130_fd_sc_hd__nor2_1
X_13024_ _03869_ _03870_ _03871_ _03786_ _03872_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__o32a_2
X_18881_ _09637_ _09675_ _09703_ VGND VGND VPWR VPWR _09773_ sky130_fd_sc_hd__o21a_1
X_10236_ net794 net60 VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__and2_1
X_17832_ _08644_ _08690_ _08641_ _08642_ VGND VGND VPWR VPWR _08693_ sky130_fd_sc_hd__nand4_2
XFILLER_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17763_ _08619_ _08620_ _08625_ VGND VGND VPWR VPWR _08626_ sky130_fd_sc_hd__o21a_1
X_14975_ _05748_ _05782_ _05869_ _05870_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__o211ai_4
X_16714_ _07435_ _07578_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__nand2_2
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17694_ _08552_ _08556_ _08555_ VGND VGND VPWR VPWR _08557_ sky130_fd_sc_hd__and3_1
X_13926_ _04696_ _04699_ _04829_ _04832_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__a31oi_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19502_ _00684_ _00686_ _00691_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_137_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16645_ _07515_ _07516_ _07512_ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__a21o_1
XFILLER_90_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19433_ _00614_ _00616_ _09199_ _09362_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13857_ _04741_ _04758_ _04729_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__a21o_1
X_16576_ _07444_ _07445_ _07447_ VGND VGND VPWR VPWR _07448_ sky130_fd_sc_hd__a21o_1
X_12808_ net659 b_h\[12\] b_h\[13\] net920 VGND VGND VPWR VPWR _03737_ sky130_fd_sc_hd__a22oi_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13788_ _04576_ _04577_ _04474_ _04691_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__a211o_1
X_19364_ _10071_ _00539_ _00540_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_33_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ net1120 net1105 VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__nand2_1
X_18315_ _09161_ _09162_ VGND VGND VPWR VPWR _09163_ sky130_fd_sc_hd__nand2_1
X_12739_ _03660_ _03662_ _03663_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__and3_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19295_ _00462_ _00453_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18246_ _09087_ _09092_ _08957_ _08958_ VGND VGND VPWR VPWR _09093_ sky130_fd_sc_hd__o2bb2ai_1
X_15458_ net640 net635 _05043_ _06312_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_100_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14409_ _05307_ _05309_ _05300_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_146_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap201 _02231_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18177_ _08962_ _08999_ _09001_ VGND VGND VPWR VPWR _09024_ sky130_fd_sc_hd__o21ai_1
X_15389_ _06237_ _06279_ _06235_ _06236_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__nand4_4
Xhold526 term_high\[62\] VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 term_low\[7\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold504 mid_sum\[29\] VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ _07989_ _07991_ _07996_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__o21ai_2
Xmax_cap234 _08230_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_2
Xmax_cap223 _06355_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
Xhold559 term_high\[56\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 term_high\[50\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap278 _07665_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_4
X_17059_ _07924_ _07927_ _07921_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__and3_1
Xmax_cap267 _03763_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_2
Xhold537 term_low\[15\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap289 _04435_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_2
X_20070_ _09308_ _09319_ _01110_ _01218_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__o22a_1
XFILLER_100_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20406_ clknet_leaf_47_clk _00046_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfxtp_1
X_20337_ net793 net32 VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__and2_2
XFILLER_107_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11070_ _02009_ net1106 net967 VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__nand3_1
XFILLER_89_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap790 net791 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__buf_12
XFILLER_115_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput68 net68 VGND VGND VPWR VPWR p[11] sky130_fd_sc_hd__buf_2
XFILLER_49_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20268_ _01479_ _01510_ _01511_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__or3_1
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput79 net79 VGND VGND VPWR VPWR p[21] sky130_fd_sc_hd__buf_2
XFILLER_102_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20199_ _01435_ net202 _01393_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__nor3_1
XFILLER_0_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _05407_ _05408_ _05532_ _05533_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__and4_1
X_11972_ net323 _02907_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__nand2_1
XFILLER_84_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13711_ _04599_ _04605_ _04614_ _04615_ _04604_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__o221a_1
XFILLER_17_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10923_ net704 net700 VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__nand2_8
X_14691_ _05583_ _05565_ _05586_ _05561_ net312 VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__o2111ai_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10854_ net793 net1263 VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__and2_1
X_16430_ _07301_ _07303_ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__nand2_1
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13642_ net289 _04486_ _04546_ _04547_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__o211ai_4
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16361_ net572 net570 net532 net528 VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__nand4_2
X_13573_ _09690_ _04481_ _04482_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__and3_1
X_10785_ p_hl\[23\] p_lh\[23\] p_hl\[22\] p_lh\[22\] VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__o211a_1
X_18100_ _08939_ _08941_ _08945_ VGND VGND VPWR VPWR _08949_ sky130_fd_sc_hd__or3_1
X_12524_ _03287_ _03290_ _03449_ net291 VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__o2bb2ai_4
X_19080_ _09966_ _09970_ VGND VGND VPWR VPWR _09971_ sky130_fd_sc_hd__nand2_1
X_15312_ _06201_ _06204_ _06202_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__a21oi_1
X_16292_ _07165_ _07166_ net281 VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__a21oi_1
X_18031_ _08868_ _08877_ _08878_ VGND VGND VPWR VPWR _08881_ sky130_fd_sc_hd__nand3_1
XFILLER_9_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12455_ _03314_ _03385_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__nand2_2
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_15243_ _06080_ _06138_ _06137_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__a21boi_1
X_11406_ _09624_ _09635_ _01855_ _02343_ _02344_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__o32ai_1
XFILLER_126_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12386_ _03310_ _03311_ _03309_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__o21ai_1
X_15174_ _06066_ _06067_ _06068_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__and3_1
XFILLER_126_777 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14125_ _05020_ _05022_ _05027_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11337_ net667 net1027 VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__nand2_8
XFILLER_141_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19982_ _01205_ _01206_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__nand2_1
XFILLER_140_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11268_ net464 _02201_ _02200_ _02199_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__o211a_1
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14056_ _04959_ _04961_ _04701_ _04818_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__o2bb2ai_4
X_18933_ _09819_ _09814_ _09810_ _09818_ VGND VGND VPWR VPWR _09825_ sky130_fd_sc_hd__o211a_1
X_11199_ _02137_ _02141_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__nand2_2
X_13007_ _03886_ _03888_ _03928_ _03930_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__o22ai_1
X_10219_ p_lh\[9\] VGND VGND VPWR VPWR _09570_ sky130_fd_sc_hd__inv_2
X_18864_ _09753_ _09754_ _09749_ VGND VGND VPWR VPWR _09756_ sky130_fd_sc_hd__a21bo_1
X_17815_ net555 net480 VGND VGND VPWR VPWR _08676_ sky130_fd_sc_hd__nand2_2
X_18795_ net606 net747 _09684_ _09685_ VGND VGND VPWR VPWR _09687_ sky130_fd_sc_hd__a22o_1
XFILLER_94_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17746_ _08471_ _08473_ _08607_ _08608_ VGND VGND VPWR VPWR _08609_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_38_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14958_ _05854_ _05856_ VGND VGND VPWR VPWR _05857_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17677_ _08449_ _08465_ _08539_ _08540_ VGND VGND VPWR VPWR _08541_ sky130_fd_sc_hd__o211ai_2
XFILLER_63_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13909_ _04811_ _04813_ _04673_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__nand3_1
X_14889_ _09384_ _09428_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__nor2_1
XFILLER_35_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16628_ _07353_ _07498_ net950 net502 _07497_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_102_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19416_ _00596_ _00597_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__nand2_1
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16559_ _07428_ _07430_ _07431_ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__nand3b_1
X_19347_ _00522_ _00523_ _00492_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_135_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19278_ _10040_ _10161_ _10177_ _10178_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__nand4_1
X_18229_ net372 _09073_ _09053_ _09056_ _09074_ VGND VGND VPWR VPWR _09076_ sky130_fd_sc_hd__o221ai_4
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold378 p_hh_pipe\[3\] VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 p_hh\[5\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold356 p_ll\[4\] VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20122_ _01292_ net331 _01306_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__o21ai_2
Xhold389 term_low\[9\] VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20053_ net568 net1013 net728 net1096 VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__and4_1
XFILLER_86_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10570_ net794 net1215 VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_24_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12240_ _02986_ _02990_ _02987_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__a21o_1
X_12171_ _02968_ _03102_ _03103_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__nand3_2
XFILLER_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11122_ net967 net525 net1052 net691 VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__a22oi_2
XFILLER_1_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15930_ _06806_ _06807_ _06789_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__a21oi_2
X_11053_ _01975_ _01980_ _01979_ _01986_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__a2bb2oi_2
X_15861_ _06651_ _06736_ _06737_ _06738_ _09690_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__o311a_1
XFILLER_103_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17600_ _08458_ _08462_ _08464_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__a21oi_1
X_14812_ _05711_ net690 net720 _05710_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__nand4_4
XFILLER_36_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15792_ _06667_ _06578_ _06664_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__nand3_1
X_18580_ net606 net1001 VGND VGND VPWR VPWR _09452_ sky130_fd_sc_hd__nand2_1
XFILLER_57_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _02885_ _02890_ _02889_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_86_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ net560 net498 net494 net565 VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__a22oi_4
X_14743_ _05463_ _05550_ _05639_ _05640_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__a22oi_1
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10906_ _09526_ _09581_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__nor2_1
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17462_ _08324_ _08326_ _08327_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__a21oi_4
X_14674_ net756 net750 net655 net649 VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__nand4_4
X_16413_ _07221_ _07286_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__nand2_2
X_11886_ _02803_ _02697_ net968 VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a21boi_2
X_13625_ _04528_ _04531_ _04532_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__nand3_4
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19201_ _10096_ _10090_ _09885_ net927 _10097_ VGND VGND VPWR VPWR _10098_ sky130_fd_sc_hd__o2111ai_4
X_17393_ _08259_ _08244_ _08240_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10837_ _01847_ _01853_ _01851_ _01852_ net795 VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__o221a_1
XFILLER_60_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19132_ _10017_ _10019_ _10013_ VGND VGND VPWR VPWR _10023_ sky130_fd_sc_hd__a21o_1
X_16344_ _07212_ _07214_ _07215_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__a21o_1
X_10768_ _01792_ _01793_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__nor2_1
X_13556_ _04463_ _04395_ net1133 VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__and3_1
XFILLER_13_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16275_ _07138_ _07147_ _07145_ net280 _07127_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_117_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12507_ _03281_ _03426_ _03437_ _03438_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__o211ai_2
X_13487_ _04333_ _04366_ _04364_ VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__a21o_1
X_19063_ _09947_ _09948_ _09937_ _09938_ VGND VGND VPWR VPWR _09954_ sky130_fd_sc_hd__o211ai_1
X_12438_ _03369_ _03370_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__and2_1
X_18014_ _09166_ _09220_ _08862_ VGND VGND VPWR VPWR _08864_ sky130_fd_sc_hd__o21ai_2
X_10699_ p_hl\[12\] p_lh\[12\] VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__nor2_1
X_15226_ _06118_ _06119_ _06121_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__a21o_1
XFILLER_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12369_ net687 net682 net483 net481 VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__nand4_1
X_15157_ _05998_ _06048_ _05997_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__a21oi_1
X_19965_ _01097_ _01157_ _01158_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__a21boi_1
X_14108_ _04925_ _05012_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__nand2_2
X_15088_ _05890_ _05881_ _05882_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18916_ _09802_ _09803_ VGND VGND VPWR VPWR _09808_ sky130_fd_sc_hd__nand2_1
X_14039_ _04944_ _04871_ _04943_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__nand3_4
XFILLER_122_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19896_ _01112_ _01114_ _01109_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__a21bo_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18847_ _09736_ _09738_ VGND VGND VPWR VPWR _09739_ sky130_fd_sc_hd__nor2_4
XFILLER_95_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18778_ _09663_ _09664_ _09654_ VGND VGND VPWR VPWR _09669_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_50_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17729_ _08518_ _08479_ _08517_ _08588_ _08589_ VGND VGND VPWR VPWR _08592_ sky130_fd_sc_hd__a32o_1
X_20740_ clknet_leaf_41_clk _00380_ VGND VGND VPWR VPWR p_ll\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20671_ clknet_leaf_5_clk _00311_ VGND VGND VPWR VPWR p_hl\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20105_ _01195_ _01196_ _01338_ _01339_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__nand4_1
X_20036_ net1073 _01263_ net203 VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__nand3_1
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_1_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _02673_ _02674_ _02572_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11671_ net646 net537 VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__nand2_1
XFILLER_41_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ net757 net751 net1076 net705 VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_40_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ net794 net1248 VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__and2_1
X_14390_ _05276_ _05278_ _05290_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_40_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10553_ net793 net1270 VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__and2_1
XFILLER_128_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13341_ _04204_ _04208_ _04250_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a21o_1
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16060_ _06934_ _06936_ _06746_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__a21o_1
Xrebuffer250 _02916_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlymetal6s2s_1
X_10484_ _01644_ _01643_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__and2b_1
XFILLER_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13272_ a_h\[0\] net763 _04181_ _04185_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__a22o_1
Xrebuffer283 _00561_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlymetal6s2s_1
X_15011_ net745 net642 _05907_ _05908_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__a22o_1
X_12223_ _03156_ _03147_ _03155_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__nand3_4
Xrebuffer294 net744 VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__buf_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12154_ net1035 _03085_ _03086_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_112_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_830 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11105_ net249 VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__inv_2
XFILLER_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19750_ _00865_ _00866_ _00953_ _00955_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__nand4_1
X_16962_ _07830_ _07831_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__nand2_1
X_12085_ _03002_ _03003_ _03013_ _03015_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__nand4_1
X_18701_ _09580_ _09583_ _09437_ VGND VGND VPWR VPWR _09585_ sky130_fd_sc_hd__a21boi_1
X_15913_ net628 net502 VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__and2_1
X_11036_ _01943_ _01974_ _01976_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__nand3_1
X_16893_ _07760_ _07762_ VGND VGND VPWR VPWR _07763_ sky130_fd_sc_hd__nand2_1
XFILLER_76_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19681_ _00876_ _00879_ _00734_ _00878_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__o211a_1
X_15844_ _06713_ _06718_ _06721_ net385 VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__o211ai_2
X_18632_ _09503_ net370 net301 _09496_ VGND VGND VPWR VPWR _09509_ sky130_fd_sc_hd__o211ai_2
X_15775_ _06584_ _06624_ _06620_ _06625_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18563_ _09423_ _09429_ _09223_ _09431_ VGND VGND VPWR VPWR _09434_ sky130_fd_sc_hd__o211ai_2
XFILLER_52_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17514_ _08210_ _08286_ _08377_ _08378_ _08290_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__o221a_1
X_12987_ net395 _03910_ _03912_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__a21o_1
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14726_ _05606_ _05607_ _05622_ _05625_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__nand4_1
X_11938_ _02649_ _02705_ _02704_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18494_ net1131 net589 VGND VGND VPWR VPWR _09358_ sky130_fd_sc_hd__nand2_1
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11869_ _02803_ _02804_ _02697_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__nand3_1
X_17445_ _08310_ net488 net578 VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__nand3_1
X_14657_ net761 net642 _05553_ _05554_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__a211oi_1
X_17376_ _08198_ _08242_ _08084_ _08136_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__a2bb2oi_1
X_13608_ net777 net673 VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__and2_1
X_14588_ _05486_ _05487_ _05476_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__a21o_1
X_16327_ net620 net815 net496 net491 _07190_ VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__a41o_1
XFILLER_119_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13539_ _09220_ _09406_ _04338_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__o21ai_1
X_19115_ _10004_ _10002_ VGND VGND VPWR VPWR _10005_ sky130_fd_sc_hd__nand2_1
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19046_ _09934_ _09927_ _09933_ VGND VGND VPWR VPWR _09937_ sky130_fd_sc_hd__nand3_4
X_16258_ _07130_ _07132_ net1090 net502 VGND VGND VPWR VPWR _07133_ sky130_fd_sc_hd__nand4_2
X_16189_ _06967_ _07063_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__nor2_1
X_15209_ _06023_ _06029_ _06100_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nand3_4
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19948_ _01166_ _01168_ _01170_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__a21o_1
X_19879_ _01094_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20723_ clknet_leaf_23_clk _00363_ VGND VGND VPWR VPWR p_lh\[25\] sky130_fd_sc_hd__dfxtp_1
X_20654_ clknet_leaf_12_clk _00294_ VGND VGND VPWR VPWR p_hh\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20585_ clknet_leaf_16_clk _00225_ VGND VGND VPWR VPWR p_hh_pipe\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12910_ _03836_ _03837_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__nand2_1
X_13890_ _04778_ _04793_ _04794_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__nand3_2
X_20019_ _01242_ _01244_ _01245_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__nand3_2
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12841_ _03762_ net267 _03765_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_100_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15560_ _06439_ _06442_ _06437_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__and3_1
X_12772_ _03611_ _03698_ _03699_ VGND VGND VPWR VPWR _03702_ sky130_fd_sc_hd__nand3_2
X_11723_ _02657_ _02658_ _02525_ _02529_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__o211a_1
X_15491_ _06380_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__inv_2
XFILLER_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14511_ _05180_ _05324_ _05372_ _05329_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_120_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11654_ net712 net983 net463 _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__a31oi_2
X_17230_ net450 _08096_ _08094_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__o21bai_4
XFILLER_42_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14442_ net736 net685 net677 net740 VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__a22oi_2
X_17161_ _08028_ _08022_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__nand2_1
X_10605_ net794 net1251 VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__and2_1
XFILLER_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11585_ net681 net507 VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__nand2_2
X_16112_ _09286_ _09581_ _06983_ _06986_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__o211ai_4
X_14373_ _09220_ _09493_ _02613_ net805 _05274_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__o221a_1
X_10536_ net795 net1292 VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__and2_1
Xmax_cap608 a_l\[5\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_12
X_17092_ _02338_ _06985_ net594 net488 _07954_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__o2111ai_4
X_13324_ net766 net705 net701 net772 VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__a22oi_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10467_ _01625_ _01626_ _01627_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__nor3_1
X_16043_ _06894_ _06916_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13255_ _04166_ _04167_ _04160_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__a21o_1
Xmax_cap619 net798 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__buf_6
X_12206_ _02864_ _02976_ _02979_ _02975_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_94_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10398_ _01565_ _01570_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__or2_1
XFILLER_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13186_ _04071_ net225 _04080_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__o21a_1
X_19802_ net574 b_l\[11\] VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__and2_1
X_12137_ _02832_ _02839_ _02840_ net399 _02843_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__a32o_2
X_17994_ _08837_ _08838_ _08840_ _08836_ VGND VGND VPWR VPWR _08845_ sky130_fd_sc_hd__o31ai_2
X_16945_ _07640_ _07643_ net977 _07813_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__o211ai_4
X_12068_ _02895_ _02897_ _02900_ _03000_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__o211ai_4
X_19733_ _00790_ _00792_ _00808_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__o21a_1
X_11019_ _01961_ _01963_ _01958_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__a21oi_2
XFILLER_64_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19664_ _00863_ _00864_ net603 net717 VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_125_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16876_ _07742_ _07744_ VGND VGND VPWR VPWR _07746_ sky130_fd_sc_hd__nor2_1
X_18615_ _09371_ _09481_ net780 net577 _09480_ VGND VGND VPWR VPWR _09490_ sky130_fd_sc_hd__o2111ai_4
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _06689_ _06691_ _06700_ _06702_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19595_ net603 net718 _00788_ _00789_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__a22oi_4
X_15758_ _06509_ _06634_ _06636_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nand3_1
X_18546_ _09118_ _09123_ _09283_ _09281_ VGND VGND VPWR VPWR _09415_ sky130_fd_sc_hd__a31o_2
X_15689_ _06455_ _06497_ _06498_ _06566_ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__nand4b_2
X_18477_ _09188_ _09264_ net457 _06605_ _09334_ VGND VGND VPWR VPWR _09339_ sky130_fd_sc_hd__o221ai_2
X_14709_ _05480_ _05609_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__nand2_1
X_17428_ _08289_ _08291_ _08290_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__nand3_2
X_17359_ _08225_ _08224_ VGND VGND VPWR VPWR _08226_ sky130_fd_sc_hd__nand2_1
XFILLER_118_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20370_ clknet_leaf_53_clk _00010_ VGND VGND VPWR VPWR b_l\[10\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_31_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload40 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__inv_8
Xclkload51 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__bufinv_16
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19029_ _09776_ _09780_ _09779_ VGND VGND VPWR VPWR _09920_ sky130_fd_sc_hd__a21boi_2
XFILLER_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ clknet_leaf_36_clk _00346_ VGND VGND VPWR VPWR p_lh\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_8_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20637_ clknet_leaf_26_clk _00277_ VGND VGND VPWR VPWR p_hh\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire138 _04090_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_8
X_11370_ _02266_ _02267_ _02309_ _02310_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__nand4_2
X_20568_ clknet_leaf_7_clk _00208_ VGND VGND VPWR VPWR mid_sum\[31\] sky130_fd_sc_hd__dfxtp_1
Xwire149 _09206_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10321_ _00891_ _00902_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__nor2_1
X_20499_ clknet_leaf_17_clk _00139_ VGND VGND VPWR VPWR term_mid\[43\] sky130_fd_sc_hd__dfxtp_1
X_13040_ _03903_ _03964_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__nand2_1
X_10252_ _09690_ net1170 VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__and2_1
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10183_ a_h\[0\] VGND VGND VPWR VPWR _09177_ sky130_fd_sc_hd__clkinv_8
XFILLER_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14991_ _05886_ _05663_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__o21ai_4
X_16730_ _07455_ _07458_ _07460_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__o21a_1
XFILLER_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13942_ _01888_ _04555_ net731 net703 _04844_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__o2111ai_2
X_16661_ _07529_ _07523_ VGND VGND VPWR VPWR _07533_ sky130_fd_sc_hd__nand2_1
XFILLER_62_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13873_ net734 net703 VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__nand2_1
X_16592_ _09199_ _09646_ _07459_ _07460_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__o211ai_1
X_15612_ _06482_ _06488_ _06490_ _06472_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o211ai_1
X_18400_ _09250_ _09251_ net604 net764 VGND VGND VPWR VPWR _09256_ sky130_fd_sc_hd__nand4_2
X_12824_ net1015 net490 _03748_ _03749_ VGND VGND VPWR VPWR _03753_ sky130_fd_sc_hd__a22o_1
XFILLER_62_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19380_ _10118_ _10134_ _00556_ _00557_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__nand4_4
X_15543_ _06423_ _06424_ _06406_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__a21oi_1
X_18331_ _09045_ _09082_ _09083_ VGND VGND VPWR VPWR _09181_ sky130_fd_sc_hd__a21boi_1
X_12755_ _03665_ _03669_ _03683_ VGND VGND VPWR VPWR _03685_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_120_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _02639_ _02605_ _02640_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__nand3_4
X_18262_ _09100_ _09101_ _09107_ VGND VGND VPWR VPWR _09109_ sky130_fd_sc_hd__a21oi_2
X_12686_ _03395_ _03407_ _03562_ _03535_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a22oi_1
X_15474_ _06346_ _06363_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__xor2_2
X_11637_ _02535_ _02531_ _02533_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__o21ai_2
X_17213_ _07936_ _07941_ _07916_ VGND VGND VPWR VPWR _08081_ sky130_fd_sc_hd__o21ai_1
X_18193_ net1128 net630 net458 _09037_ _09038_ VGND VGND VPWR VPWR _09040_ sky130_fd_sc_hd__a32o_1
X_14425_ _05321_ _05323_ _05181_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__a21oi_1
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17144_ _07857_ net472 net844 _07855_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_96_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ _09482_ _09592_ _02501_ _02503_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__o211ai_1
X_14356_ _05258_ _05259_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__nor2_1
XFILLER_7_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10519_ net1321 net1352 VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__nand2_1
XFILLER_128_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap405 _01812_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
X_17075_ _07936_ _07938_ _07917_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__o21ai_1
Xmax_cap416 _08375_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_2
X_13307_ net777 net693 VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nand2_1
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11499_ _02436_ _02434_ _02433_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__and3_1
X_16026_ _06900_ _06902_ _09144_ _09613_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__o2bb2ai_1
Xmax_cap438 _02874_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__buf_1
Xmax_cap449 _08169_ VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_6
X_14287_ net703 net699 _05043_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__and3_1
XFILLER_143_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13238_ _04144_ _04153_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__xor2_1
XFILLER_111_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13169_ _03950_ _03952_ _03951_ _04091_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a31oi_4
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17977_ _08827_ _08828_ VGND VGND VPWR VPWR _08829_ sky130_fd_sc_hd__nor2_1
X_19716_ net1079 net574 net1033 net567 _00912_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__a41o_1
X_16928_ _09253_ _09613_ _07669_ _07672_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__o31a_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16859_ _07724_ _07727_ _07725_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__nand3_1
X_19647_ _00845_ _00847_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__nand2_1
XFILLER_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19578_ _00671_ _00673_ _00643_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_105_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18529_ _09388_ _09391_ _09350_ _09386_ VGND VGND VPWR VPWR _09397_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_47_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20422_ clknet_leaf_18_clk net139 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20353_ net794 net50 VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__and2_1
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20284_ _09362_ _09373_ _01529_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__or3_1
XFILLER_121_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10870_ net793 net1303 VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__and2_1
XFILLER_45_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12540_ _03469_ _03470_ _03465_ VGND VGND VPWR VPWR _03472_ sky130_fd_sc_hd__and3_1
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12471_ _03398_ net483 net679 net687 net475 VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__a32oi_2
X_11422_ net659 net873 VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__nand2_4
X_14210_ net714 b_l\[15\] _05109_ _05112_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__a22o_1
X_15190_ _02278_ net455 _06013_ _06040_ _06084_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_78_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14141_ net728 net724 net709 net703 VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__nand4_1
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11353_ net681 net1061 net525 net1052 VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__and4_1
X_11284_ _02216_ _02219_ _02224_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__nand3_1
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14072_ _02362_ _04182_ _04973_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__o21ai_2
X_10304_ term_low\[21\] term_mid\[21\] _00719_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__o21ai_1
X_17900_ net253 _08754_ _08757_ VGND VGND VPWR VPWR _08759_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_91_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13023_ _03791_ _03875_ _03786_ _03789_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__nand4_4
XFILLER_79_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18880_ _09677_ _09703_ VGND VGND VPWR VPWR _09772_ sky130_fd_sc_hd__nand2_1
X_10235_ net794 net59 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__and2_1
X_17831_ _08691_ VGND VGND VPWR VPWR _08692_ sky130_fd_sc_hd__inv_2
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17762_ _08622_ _08277_ _08273_ VGND VGND VPWR VPWR _08625_ sky130_fd_sc_hd__nand3_4
XFILLER_47_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14974_ _05871_ _05866_ _05872_ _05783_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__o211ai_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16713_ _07438_ _07583_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__nand2_4
XFILLER_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17693_ net1093 net476 VGND VGND VPWR VPWR _08556_ sky130_fd_sc_hd__and2_1
X_13925_ _04694_ _04829_ _04831_ _09690_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__o31ai_1
X_19501_ _00488_ _00688_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_122_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16644_ net570 net936 net947 net523 VGND VGND VPWR VPWR _07516_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_89_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13856_ _04736_ net1132 _04758_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__o21ai_2
X_19432_ _00612_ _00613_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__nand2_1
XFILLER_90_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12807_ net669 net659 b_h\[12\] net481 VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__and4_1
X_16575_ a_l\[0\] net472 VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__nand2_1
X_10999_ net707 net517 VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__nand2_1
XFILLER_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13787_ _04692_ _04693_ _04579_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__a21bo_1
X_19363_ _00534_ _10114_ _10070_ _00535_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__nand4_4
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ net797 _06409_ _06410_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__nor3_1
X_18314_ _09156_ _09157_ _09147_ VGND VGND VPWR VPWR _09162_ sky130_fd_sc_hd__nand3_2
X_12738_ net321 _03656_ _03657_ _03664_ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a31o_1
X_19294_ _00454_ _00465_ _00466_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__nand3_4
X_12669_ _03597_ _03599_ _03499_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_100_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18245_ _09090_ _09024_ _09088_ VGND VGND VPWR VPWR _09092_ sky130_fd_sc_hd__nand3_1
X_15457_ net722 net719 net640 net635 VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_100_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _05308_ _05310_ _05299_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18176_ _08894_ _08950_ _09022_ _09023_ net794 VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__o311a_1
X_15388_ _06238_ _06278_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__nand2_1
Xmax_cap202 _01437_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__buf_1
Xmax_cap213 _01990_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
Xhold505 mid_sum\[28\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
X_17127_ _07994_ _07988_ VGND VGND VPWR VPWR _07996_ sky130_fd_sc_hd__nand2_2
Xmax_cap235 _08129_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
Xhold516 p_ll\[28\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
X_14339_ _05186_ _05190_ _05233_ _05235_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__nand4_1
Xmax_cap224 _06195_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__buf_2
Xhold549 _00066_ VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap268 _03069_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
X_17058_ net571 net561 net964 net506 VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__nand4_1
Xhold538 p_ll\[29\] VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16009_ _09210_ _09602_ _06537_ _06880_ _06879_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__o221a_4
Xmax_cap279 _07663_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20405_ clknet_leaf_43_clk _00045_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20336_ net793 net31 VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__and2_2
Xmax_cap791 net792 VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__buf_12
Xmax_cap780 b_l\[2\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_73_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput69 net69 VGND VGND VPWR VPWR p[12] sky130_fd_sc_hd__buf_2
X_20267_ _01510_ _01511_ _01475_ _01478_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20198_ _01435_ net202 _01393_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11971_ _02903_ _02902_ _02892_ VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__nand3_4
XFILLER_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10922_ net697 net545 net538 net702 VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__a22o_1
XFILLER_84_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13710_ net456 _04613_ _04616_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__o21a_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14690_ _05564_ _05587_ _05588_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__nand3_1
X_10853_ net793 net1209 VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__and2_1
X_13641_ _04546_ _04547_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__nand2_2
XFILLER_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10784_ _01806_ _01807_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__or2_1
XFILLER_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16360_ net577 net569 VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__nand2_8
X_13572_ _04389_ _04477_ _04387_ _04388_ _04479_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__a221o_1
X_16291_ _07024_ _07039_ _07159_ _07158_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__o211ai_4
X_12523_ _03287_ _03290_ _03450_ _03452_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__and4_1
XFILLER_40_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15311_ _06201_ _06203_ _06204_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__a21o_1
X_18030_ _08840_ _08866_ _08875_ _08876_ VGND VGND VPWR VPWR _08880_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_9_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15242_ _06082_ _06133_ _06134_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__nand3_2
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12454_ net661 net995 net495 net665 VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a22oi_1
X_11405_ _02343_ _02344_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__nor2_1
X_12385_ _09449_ _09646_ _03310_ _03311_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__o22a_1
X_15173_ _06064_ _06065_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__nand3_1
XFILLER_126_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11336_ _02170_ _02275_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__nand2_2
X_14124_ _05019_ _05021_ _05008_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__a21oi_1
X_19981_ _09297_ _09329_ _09351_ _09286_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__o22a_1
XFILLER_141_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14055_ _04955_ _04957_ _04958_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__nand3_2
X_18932_ _09822_ _09809_ _09821_ VGND VGND VPWR VPWR _09824_ sky130_fd_sc_hd__nand3_2
XFILLER_140_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11267_ _02199_ net361 net440 VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__a21bo_1
X_13006_ _03887_ _03889_ _03929_ _03931_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__nand4_1
X_11198_ _02131_ _02134_ _02133_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__nand3_2
XFILLER_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10218_ p_hl\[9\] VGND VGND VPWR VPWR _09559_ sky130_fd_sc_hd__inv_2
X_18863_ net619 net732 _09753_ _09754_ VGND VGND VPWR VPWR _09755_ sky130_fd_sc_hd__a22oi_4
X_17814_ a_l\[12\] net477 VGND VGND VPWR VPWR _08675_ sky130_fd_sc_hd__and2_1
X_18794_ _09684_ _09685_ net606 net747 VGND VGND VPWR VPWR _09686_ sky130_fd_sc_hd__nand4_1
X_17745_ _08549_ _08602_ _08603_ VGND VGND VPWR VPWR _08608_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_38_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14957_ _05714_ _05727_ _05726_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__a21boi_2
X_17676_ _08533_ _08534_ _08536_ VGND VGND VPWR VPWR _08540_ sky130_fd_sc_hd__a21o_1
XFILLER_63_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13908_ _04813_ _04673_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__nand2_1
X_14888_ _05710_ _05712_ _05733_ _05738_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__a22o_1
XFILLER_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16627_ net590 net1069 net513 net506 VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_102_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19415_ net579 net744 net738 net588 VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__a22oi_4
X_13839_ net783 net656 net650 net788 VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__a22oi_4
X_16558_ _07292_ _07294_ _07289_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__a21boi_2
XFILLER_50_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19346_ _00494_ _00520_ _00521_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__nand3_4
X_15509_ _06392_ _06395_ _06390_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_135_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16489_ _07359_ _07360_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__a21oi_1
X_19277_ _10177_ _10178_ VGND VGND VPWR VPWR _10179_ sky130_fd_sc_hd__nand2_1
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18228_ net372 _09073_ _09074_ VGND VGND VPWR VPWR _09075_ sky130_fd_sc_hd__o21ai_2
XFILLER_116_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18159_ _08963_ _08997_ _08998_ net337 VGND VGND VPWR VPWR _09007_ sky130_fd_sc_hd__a31o_1
Xhold368 p_ll_pipe\[6\] VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 term_low\[3\] VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20121_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__inv_2
XFILLER_131_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold379 p_ll_pipe\[24\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_86_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20052_ net563 net724 VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__nand2_1
XFILLER_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12170_ _02968_ _03103_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__nand2_1
XFILLER_108_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11121_ net686 net525 VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__nand2_1
XFILLER_122_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20319_ net793 net16 VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__and2_1
X_11052_ _01986_ _01979_ _01975_ _01980_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15860_ _06651_ _06737_ _06736_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__o21ai_1
XFILLER_103_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14811_ _05604_ _05709_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nand2_1
X_15791_ _06664_ _06667_ _06505_ _06577_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11954_ _02883_ _02888_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__nand2_2
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ net560 net500 VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__nand2_2
X_14742_ _05463_ _05550_ _05639_ _05640_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__nand4_2
X_11885_ _02797_ _02798_ _02802_ _02804_ _02698_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a32oi_2
X_17461_ _08205_ _08220_ _08218_ _08214_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__o2bb2ai_4
X_10905_ a_h\[0\] net1076 VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__nand2_4
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14673_ net750 net756 net655 net649 VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__and4_1
X_16412_ net257 net256 _07283_ VGND VGND VPWR VPWR _07286_ sky130_fd_sc_hd__nand3_4
X_10836_ _01849_ _01850_ p_hl\[30\] p_lh\[30\] VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_72_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13624_ _04415_ _04526_ _04523_ _04517_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__a22oi_2
XFILLER_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19200_ _10089_ _10091_ _09210_ _09308_ VGND VGND VPWR VPWR _10097_ sky130_fd_sc_hd__o2bb2ai_1
X_17392_ _08249_ _08253_ _08256_ VGND VGND VPWR VPWR _08259_ sky130_fd_sc_hd__o21ai_1
X_19131_ _10017_ _10019_ _09253_ _09264_ VGND VGND VPWR VPWR _10022_ sky130_fd_sc_hd__o2bb2ai_1
X_16343_ _07212_ _07214_ _07215_ VGND VGND VPWR VPWR _07217_ sky130_fd_sc_hd__a21oi_1
X_10767_ p_hl\[22\] p_lh\[22\] VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__nor2_1
X_13555_ net1133 _04463_ _04395_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16274_ _07138_ _07147_ _07145_ VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_117_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12506_ _03434_ _03428_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__nand2_1
X_13486_ _04395_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__inv_2
X_10698_ _09690_ _01733_ _01734_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__and3_1
X_19062_ _09947_ _09948_ _09937_ _09938_ VGND VGND VPWR VPWR _09953_ sky130_fd_sc_hd__o211a_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12437_ _03362_ _03367_ _03364_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__nand3_1
X_18013_ _04182_ _06441_ net630 net764 _08861_ VGND VGND VPWR VPWR _08863_ sky130_fd_sc_hd__o2111ai_4
XFILLER_9_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15225_ _06030_ _06026_ _06015_ _06032_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__o22a_2
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15156_ _06050_ _06051_ _05997_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_130_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12368_ net687 net682 net483 net481 VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__and4_1
X_14107_ net756 net670 VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__nand2_2
X_12299_ _03218_ _03219_ _03230_ VGND VGND VPWR VPWR _03233_ sky130_fd_sc_hd__a21o_1
X_11319_ _02190_ _02255_ net706 net501 _02258_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__o2111ai_1
XFILLER_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19964_ _01094_ _01096_ _01157_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__a21boi_2
X_15087_ _05982_ _05984_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__nand2_1
XFILLER_141_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18915_ net446 _09806_ _09804_ VGND VGND VPWR VPWR _09807_ sky130_fd_sc_hd__o21ai_1
X_19895_ _01020_ _01110_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__nand2_1
X_14038_ _04913_ _04916_ _04936_ net317 VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18846_ _09329_ _09351_ _06402_ _09626_ _09630_ VGND VGND VPWR VPWR _09738_ sky130_fd_sc_hd__o311a_1
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15989_ net1116 net529 VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__nand2_1
X_18777_ _09483_ net412 _09665_ _09666_ VGND VGND VPWR VPWR _09667_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_50_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17728_ _08513_ _08516_ _08588_ _08589_ _08519_ VGND VGND VPWR VPWR _08591_ sky130_fd_sc_hd__o2111ai_2
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17659_ _08519_ _08517_ _08426_ _08521_ VGND VGND VPWR VPWR _08523_ sky130_fd_sc_hd__a211oi_1
XFILLER_63_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20670_ clknet_leaf_5_clk _00310_ VGND VGND VPWR VPWR p_hl\[4\] sky130_fd_sc_hd__dfxtp_2
X_19329_ _00501_ net732 net598 VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__nand3_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20104_ _01195_ _01196_ _01338_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__a22o_1
XFILLER_86_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20035_ _09242_ _09384_ _01092_ _01090_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__o31ai_1
XFILLER_86_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11670_ net652 net535 VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__nand2_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ clknet_leaf_2_clk _00439_ VGND VGND VPWR VPWR b_h\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ net794 net1156 VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10552_ net793 net1269 VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__and2_1
X_13340_ _04248_ _04249_ _04252_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__a21o_1
Xrebuffer240 b_h\[2\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd1_1
X_13271_ net923 net953 net710 net704 VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__nand4_1
X_10483_ _01641_ _01642_ _01636_ net796 VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__a31o_1
XFILLER_136_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12222_ _03150_ _03152_ _03148_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__a21bo_1
X_15010_ _05797_ _05906_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__nand2_1
XFILLER_123_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer284 _09677_ VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__buf_6
Xrebuffer295 net744 VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__buf_2
X_12153_ _03087_ _03083_ _03082_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_112_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_842 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11104_ _02034_ _02035_ net991 _02044_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16961_ _07655_ _07658_ _07827_ _07828_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__nand4_4
X_12084_ _03002_ net357 _03012_ _03014_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_78_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15912_ _06660_ _06788_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__nor2_1
X_11035_ _01928_ _01941_ _01954_ _01973_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18700_ _09580_ _09583_ VGND VGND VPWR VPWR _09584_ sky130_fd_sc_hd__nand2_1
X_16892_ _07759_ net452 _07748_ _07758_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__o211ai_4
X_19680_ _00881_ _00735_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__nand2_1
X_15843_ _06721_ _06720_ net386 VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__a21o_1
XFILLER_94_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18631_ _09506_ _09507_ VGND VGND VPWR VPWR _09508_ sky130_fd_sc_hd__nor2_1
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15774_ _06508_ _06634_ _06635_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__a21o_1
X_18562_ _09431_ _09223_ VGND VGND VPWR VPWR _09433_ sky130_fd_sc_hd__nand2_1
X_12986_ _03909_ _03910_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__a21oi_2
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17513_ net550 net969 net504 net554 VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__a22oi_2
X_14725_ _05606_ _05607_ _05625_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_28_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11937_ _02871_ _02869_ _02866_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__nand3_2
X_18493_ _09355_ _09356_ VGND VGND VPWR VPWR _09357_ sky130_fd_sc_hd__nand2_1
X_11868_ _02695_ _02696_ _02803_ _02804_ VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__a2bb2o_1
X_17444_ net569 net565 net498 net493 VGND VGND VPWR VPWR _08310_ sky130_fd_sc_hd__nand4_2
X_14656_ net771 net767 net640 net636 _05552_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__a41o_1
XFILLER_33_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11799_ net1036 net546 net537 net644 VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a22oi_2
X_10819_ _01832_ _01837_ _01838_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__o21a_1
X_17375_ _08200_ net234 _08232_ VGND VGND VPWR VPWR _08242_ sky130_fd_sc_hd__nand3_1
X_13607_ _04509_ _04514_ _04513_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__o21ai_2
X_14587_ _05472_ _05474_ _05486_ _05487_ VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__nand4_1
X_16326_ net841 net1032 _07194_ _07196_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19114_ _09734_ _10003_ _09733_ _09730_ VGND VGND VPWR VPWR _10004_ sky130_fd_sc_hd__nand4_4
X_13538_ _09220_ _09406_ _04338_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__o21a_1
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19045_ _09931_ _09932_ net883 net557 VGND VGND VPWR VPWR _09936_ sky130_fd_sc_hd__nand4_2
X_16257_ net607 net966 net512 net505 VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__nand4_1
X_13469_ _04258_ _04304_ _04305_ _04309_ _04214_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a32o_1
XFILLER_133_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16188_ _06956_ _06963_ _06964_ _06971_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__a31oi_4
X_15208_ _06023_ _06029_ _06100_ _06102_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__a22o_1
X_15139_ _06034_ _06015_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__nand2_1
XFILLER_99_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19947_ _01170_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__inv_2
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19878_ _01093_ net591 _01090_ net717 VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_143_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18829_ _09554_ _09556_ _09716_ _09717_ VGND VGND VPWR VPWR _09722_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_26_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20722_ clknet_leaf_23_clk _00362_ VGND VGND VPWR VPWR p_lh\[24\] sky130_fd_sc_hd__dfxtp_1
X_20653_ clknet_leaf_12_clk _00293_ VGND VGND VPWR VPWR p_hh\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire309 _06528_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_63_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20584_ clknet_leaf_16_clk _00224_ VGND VGND VPWR VPWR p_hh_pipe\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20018_ net332 _01136_ _01240_ _01105_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__a22oi_2
X_12840_ _03654_ _03764_ net267 _03762_ VGND VGND VPWR VPWR _03769_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_83_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12771_ _03612_ _03696_ _03697_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__nand3b_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11722_ _02525_ _02529_ _02657_ _02658_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__a211oi_2
XFILLER_70_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15490_ _06358_ _06360_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__nand2b_1
XFILLER_14_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14510_ _05378_ _05396_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nand2_1
X_11653_ net983 net483 net481 net712 VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a22oi_2
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14441_ net740 net677 VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__nand2_1
X_17160_ _07584_ _08024_ _07586_ _08022_ _08027_ VGND VGND VPWR VPWR _08029_ sky130_fd_sc_hd__a311o_1
XFILLER_80_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10604_ net794 net1275 VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__and2_1
X_14372_ net771 net767 net649 net642 VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__nand4_2
X_11584_ _02397_ _02522_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__nand2_1
X_16111_ _06983_ _06986_ _06980_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__a21o_1
X_13323_ net772 net766 net705 net701 VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__nand4_2
X_10535_ net795 net1171 VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__and2_1
X_17091_ _09253_ _09275_ _02338_ _07951_ _07954_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__o311a_1
Xmax_cap609 net610 VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_12
X_10466_ _01626_ _01627_ _01625_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__o21a_1
X_16042_ _06894_ _06911_ _06912_ _06916_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__nand4_1
XFILLER_129_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13254_ _04166_ _04167_ _04160_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12205_ _03127_ _03134_ _03135_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__nand3_4
X_13185_ _04105_ _04106_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__nand2_1
X_10397_ net167 _01566_ _01569_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__o21ai_2
X_12136_ _02831_ _02843_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__and2_1
X_19801_ _00919_ _00911_ _00917_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__a21boi_1
X_17993_ _09144_ _09155_ _08838_ _08840_ VGND VGND VPWR VPWR _08844_ sky130_fd_sc_hd__o22a_1
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16944_ _07640_ _07643_ _07813_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__o21ai_2
X_12067_ _02898_ _02904_ _02997_ _02998_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__nand4_4
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19732_ _00934_ _00897_ _00933_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__nand3_4
X_11018_ net967 net681 net965 net538 VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nand4_4
X_16875_ net798 net476 _07740_ _07741_ VGND VGND VPWR VPWR _07745_ sky130_fd_sc_hd__a22o_1
X_19663_ net603 net717 _00863_ _00864_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__a22o_1
XFILLER_37_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _06689_ _06691_ _06701_ _06703_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__nand4_1
XFILLER_92_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18614_ _09297_ _09319_ net459 _09480_ _09486_ VGND VGND VPWR VPWR _09489_ sky130_fd_sc_hd__o311a_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19594_ _09210_ _09362_ _00787_ _00789_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__or4b_1
X_15757_ _06634_ _06636_ VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__nand2_1
XFILLER_92_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18545_ _09412_ _09413_ VGND VGND VPWR VPWR _09414_ sky130_fd_sc_hd__nand2_2
X_12969_ _03895_ _03890_ _03892_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__and3_1
X_15688_ _06560_ _06563_ _06455_ _06499_ VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__a211oi_1
X_18476_ net619 net1148 _09334_ _09335_ VGND VGND VPWR VPWR _09338_ sky130_fd_sc_hd__a22o_1
X_14708_ _05478_ _05481_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__nand2_1
X_17427_ _08289_ _08291_ _08290_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__and3_1
X_14639_ _05517_ _05507_ _05506_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__a21boi_2
XFILLER_21_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17358_ _08217_ _08205_ _08041_ VGND VGND VPWR VPWR _08225_ sky130_fd_sc_hd__a21oi_1
X_16309_ _07060_ _07181_ _07182_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__and3_1
X_17289_ _08149_ _08148_ _08010_ _08155_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_31_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload52 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__bufinv_16
Xclkload41 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__inv_6
XFILLER_115_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload30 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_6
X_19028_ _09917_ _09918_ VGND VGND VPWR VPWR _09919_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20705_ clknet_leaf_34_clk _00345_ VGND VGND VPWR VPWR p_lh\[7\] sky130_fd_sc_hd__dfxtp_1
Xwire139 _00062_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
X_20636_ clknet_leaf_26_clk _00276_ VGND VGND VPWR VPWR p_hh\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload2 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
X_20567_ clknet_leaf_7_clk _00207_ VGND VGND VPWR VPWR mid_sum\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10320_ term_low\[25\] term_mid\[25\] VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__and2_1
X_20498_ clknet_leaf_17_clk _00138_ VGND VGND VPWR VPWR term_mid\[42\] sky130_fd_sc_hd__dfxtp_1
X_10251_ _09690_ net1199 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10182_ net974 VGND VGND VPWR VPWR _09166_ sky130_fd_sc_hd__clkinv_8
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14990_ _05664_ _05886_ _05885_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__o21a_4
X_13941_ _04844_ _04845_ _09308_ _09395_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_115_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16660_ _07527_ net970 net876 net541 VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__nand4_2
X_13872_ net731 net709 VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__nand2_2
XFILLER_35_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16591_ _07459_ _07460_ _07455_ VGND VGND VPWR VPWR _07463_ sky130_fd_sc_hd__a21o_1
X_15611_ _06448_ _06461_ _06491_ _06492_ VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__o211ai_2
XFILLER_74_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12823_ _03748_ _03749_ net1015 net490 VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__nand4_1
XFILLER_62_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15542_ net1062 _06402_ _06408_ _06425_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__or4b_1
X_18330_ _09081_ _09080_ _09078_ _09083_ net277 VGND VGND VPWR VPWR _09180_ sky130_fd_sc_hd__a32oi_4
X_12754_ _03661_ _03668_ _03682_ _03666_ VGND VGND VPWR VPWR _03684_ sky130_fd_sc_hd__o211ai_2
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ net325 _02624_ _02631_ _02634_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o2bb2ai_4
X_18261_ _09105_ _09102_ _09106_ VGND VGND VPWR VPWR _09108_ sky130_fd_sc_hd__o21a_1
X_17212_ _07912_ _07898_ _07939_ _07937_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__o211ai_1
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12685_ _03397_ _03550_ _03554_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__o21ai_2
X_15473_ _06346_ _06363_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__and2b_1
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11636_ _09177_ _09657_ _02462_ _02461_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__o31ai_1
X_18192_ net458 _06401_ _09037_ _09038_ VGND VGND VPWR VPWR _09039_ sky130_fd_sc_hd__a22oi_1
X_14424_ _05297_ _05298_ _05316_ _05317_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__o2bb2ai_1
X_17143_ _08009_ _08011_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__nand2_1
X_11567_ _09526_ _09581_ _02502_ _02501_ _02497_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_96_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _05100_ _05105_ _05257_ net796 VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__a31o_1
X_10518_ net1372 _01660_ _01664_ net1352 VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__a31o_1
X_17074_ _07917_ _07937_ _07939_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__nand3_1
X_13306_ _04192_ _04197_ _04193_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__a21oi_1
Xmax_cap406 _00764_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_2
X_14286_ _05034_ _05187_ _05188_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__nand3_4
X_11498_ _02433_ _02434_ _02436_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__a21oi_4
X_16025_ net1127 net613 net512 net505 VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__nand4_2
Xmax_cap439 _02299_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
X_13237_ _04151_ _04152_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__nand2b_1
XFILLER_6_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10449_ term_mid\[43\] term_high\[43\] term_mid\[42\] term_high\[42\] VGND VGND VPWR
+ VPWR _01614_ sky130_fd_sc_hd__o211a_1
XFILLER_130_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13168_ _03944_ _03947_ _04089_ _03948_ _03997_ VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__o2111ai_1
X_12119_ net679 net492 VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__nand2_1
X_17976_ _08825_ _08826_ net632 net774 VGND VGND VPWR VPWR _08828_ sky130_fd_sc_hd__and4_1
X_13099_ _03983_ _04023_ _03984_ _03976_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__nand4_2
X_16927_ net376 _07795_ _07790_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__o21ai_1
X_19715_ _09275_ _09308_ _00920_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__o21ai_2
XFILLER_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16858_ _07724_ _07727_ VGND VGND VPWR VPWR _07729_ sky130_fd_sc_hd__nand2_1
XFILLER_93_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19646_ _00584_ _00587_ _00843_ _00844_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__o211ai_2
X_15809_ _06680_ _06683_ _06677_ VGND VGND VPWR VPWR _06688_ sky130_fd_sc_hd__a21o_1
X_16789_ net378 _07654_ _07636_ net344 VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__o211ai_2
XFILLER_1_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19577_ _00770_ _00771_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18528_ _09393_ _09350_ VGND VGND VPWR VPWR _09396_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_47_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18459_ _09316_ _09320_ net797 VGND VGND VPWR VPWR _09321_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_16_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20421_ clknet_leaf_27_clk _00061_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20352_ net794 net49 VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__and2_1
XFILLER_134_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20283_ net716 _01410_ _01528_ net724 VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__o22a_1
XFILLER_114_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12470_ _03300_ _03397_ net687 net475 _03400_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__o2111a_1
XFILLER_8_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11421_ _02358_ _02359_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__nand2_2
X_20619_ clknet_leaf_42_clk _00259_ VGND VGND VPWR VPWR p_ll_pipe\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11352_ net678 net525 VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14140_ net728 net724 net709 net703 VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__and4_1
X_10303_ _00536_ _00569_ _00633_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__nand3_1
X_11283_ _02224_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14071_ net771 net767 net662 net656 VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nand4_1
XFILLER_106_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13022_ _03944_ _03947_ _03948_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_5_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10234_ net794 net58 VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__and2_1
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17830_ _08645_ _08689_ VGND VGND VPWR VPWR _08691_ sky130_fd_sc_hd__nand2_1
XFILLER_79_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17761_ _07587_ _08276_ _08623_ VGND VGND VPWR VPWR _08624_ sky130_fd_sc_hd__a21oi_4
XFILLER_47_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14973_ _05867_ _05868_ _05791_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__a21o_1
X_19500_ _00488_ _00530_ _00531_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__nand3_2
X_16712_ _07582_ _07577_ net145 VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__a21oi_4
X_17692_ a_l\[11\] net565 net485 net479 VGND VGND VPWR VPWR _08555_ sky130_fd_sc_hd__nand4_1
X_13924_ _04485_ _04580_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_122_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16643_ _06999_ _07513_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13855_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__inv_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19431_ _09231_ _09329_ _09351_ _09210_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__o22a_1
X_12806_ _03734_ VGND VGND VPWR VPWR _03735_ sky130_fd_sc_hd__inv_2
X_19362_ _00538_ _00539_ _00540_ _10071_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__a22oi_1
X_16574_ _07444_ _07445_ VGND VGND VPWR VPWR _07446_ sky130_fd_sc_hd__nand2_1
X_10998_ _01915_ _01923_ net404 _01927_ _01914_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__a32o_1
XFILLER_90_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18313_ _09065_ _09146_ _09158_ _09159_ VGND VGND VPWR VPWR _09161_ sky130_fd_sc_hd__o211ai_2
X_13786_ _04475_ _04574_ _04575_ _04692_ _04693_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__a32oi_4
XFILLER_31_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _06407_ _01856_ _06406_ _06401_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__and4_1
X_12737_ net321 _03656_ _03657_ _03664_ VGND VGND VPWR VPWR _03667_ sky130_fd_sc_hd__a31oi_2
X_19293_ _09264_ _09275_ _00458_ _00460_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__o211ai_2
XFILLER_31_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12668_ _03588_ _03595_ _03598_ VGND VGND VPWR VPWR _03599_ sky130_fd_sc_hd__o21ai_1
X_18244_ _09000_ _09007_ _09088_ VGND VGND VPWR VPWR _09091_ sky130_fd_sc_hd__nand3_2
X_15456_ net719 net640 net635 net722 VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__a22oi_1
X_11619_ _02553_ _02554_ _02352_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_100_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18175_ _08894_ _08950_ _09020_ _09021_ VGND VGND VPWR VPWR _09023_ sky130_fd_sc_hd__a2bb2o_1
X_14407_ _09264_ _09460_ _09482_ _05304_ _05303_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__o221ai_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17126_ _07947_ _07986_ _07987_ _07990_ VGND VGND VPWR VPWR _07995_ sky130_fd_sc_hd__nand4_2
X_12599_ _03526_ _03529_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__nand2_1
X_15387_ _09504_ _09515_ net455 _06225_ _06238_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__o311a_1
Xhold517 p_ll_pipe\[8\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold506 p_hh\[30\] VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap225 _04081_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_1
X_14338_ _05119_ _05238_ net194 VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nand3_2
XFILLER_144_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap258 _07087_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_133_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap269 _02354_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
Xmax_cap247 _02941_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__buf_4
Xmax_cap236 _07693_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_2
Xhold528 mid_sum\[30\] VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ net571 net561 net964 net506 VGND VGND VPWR VPWR _07926_ sky130_fd_sc_hd__and4_1
X_14269_ _05155_ _05168_ _05170_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__nand3_2
Xhold539 mid_sum\[12\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16008_ _06882_ _06879_ _09210_ _09602_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__a211oi_2
XFILLER_124_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17959_ net627 net632 _04133_ _08812_ net797 VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__a311oi_1
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19629_ _00777_ _00779_ _00823_ _00826_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__a22oi_1
XFILLER_53_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_8
X_20404_ clknet_leaf_43_clk _00044_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfxtp_1
X_20335_ net793 net30 VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap781 net782 VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__buf_12
Xmax_cap770 b_l\[4\] VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__buf_12
X_20266_ _01506_ _01507_ _01508_ _01509_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__and4bb_1
XFILLER_102_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap792 b_l\[0\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__buf_12
X_20197_ _01435_ net202 _01393_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__o21a_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11970_ _02904_ _02897_ _02893_ _02905_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__o211ai_2
X_10921_ net697 net545 net538 net702 VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__a22oi_1
XFILLER_57_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10852_ net793 net1238 VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__and2_1
XFILLER_72_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13640_ _04503_ _04545_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__nand2_1
X_10783_ net1349 p_lh\[24\] VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__nor2_1
X_13571_ _04387_ _04388_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__nand3_1
X_16290_ _07163_ _07062_ _07162_ VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__nand3_4
X_12522_ _03286_ _03158_ _03452_ _03290_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o211ai_2
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_8
X_15310_ _06201_ _06203_ _06204_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__nand3_1
X_15241_ _06049_ net174 _06129_ _06135_ _06136_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__o221ai_4
X_12453_ net661 net995 VGND VGND VPWR VPWR _03385_ sky130_fd_sc_hd__nand2_1
X_11404_ _02341_ net1032 net712 _02340_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__and4b_1
X_12384_ _03315_ net489 net679 VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__nand3_1
X_15172_ _05975_ _05979_ _05976_ _05971_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__o2bb2ai_1
X_11335_ net658 net965 net539 net664 VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a22oi_4
X_19980_ net574 net1095 VGND VGND VPWR VPWR _01206_ sky130_fd_sc_hd__nand2_1
X_14123_ _05019_ _05021_ _05007_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__and3_1
XFILLER_137_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11266_ _02108_ _02109_ _02199_ net361 net464 VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__a221oi_1
XFILLER_98_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14054_ _04955_ _04957_ _04958_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__and3_1
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18931_ _09822_ _09809_ VGND VGND VPWR VPWR _09823_ sky130_fd_sc_hd__nand2_1
X_10217_ p_lh\[6\] VGND VGND VPWR VPWR _09548_ sky130_fd_sc_hd__inv_2
X_13005_ _03856_ _03927_ _03889_ _03887_ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__o211ai_1
X_11197_ _02132_ _02128_ _02054_ _02052_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__a22oi_2
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18862_ net609 net603 net1091 net737 VGND VGND VPWR VPWR _09754_ sky130_fd_sc_hd__nand4_4
XFILLER_95_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17813_ _08494_ net490 a_l\[15\] VGND VGND VPWR VPWR _08674_ sky130_fd_sc_hd__and3_1
X_18793_ net597 net760 net596 net1001 VGND VGND VPWR VPWR _09685_ sky130_fd_sc_hd__nand4_4
X_17744_ _08548_ _08604_ _08606_ VGND VGND VPWR VPWR _08607_ sky130_fd_sc_hd__nand3_1
XFILLER_48_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14956_ _05714_ _05727_ _05726_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit289 b_l\[1\] VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_38_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13907_ _04811_ _04813_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__nand2_1
XFILLER_48_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17675_ _08533_ _08534_ _08536_ VGND VGND VPWR VPWR _08539_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_59_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14887_ _05710_ _05712_ _05733_ _05738_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__a22oi_1
X_19414_ net579 net835 VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__nand2_1
X_16626_ net584 net506 VGND VGND VPWR VPWR _07498_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_102_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13838_ net788 net650 VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__nand2_1
X_16557_ _07421_ _07423_ _07427_ VGND VGND VPWR VPWR _07430_ sky130_fd_sc_hd__nand3_1
X_13769_ _04670_ _04671_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_44_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19345_ _00505_ _00518_ _00507_ _00516_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__o211ai_2
Xclkbuf_leaf_42_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_8
X_15508_ _06392_ _06395_ _06390_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__o21a_1
X_19276_ _09373_ _10163_ _10173_ _10174_ VGND VGND VPWR VPWR _10178_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_135_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16488_ _07246_ _07242_ _07245_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__o21ai_2
X_18227_ _09069_ _09070_ _09060_ VGND VGND VPWR VPWR _09074_ sky130_fd_sc_hd__nand3_4
X_15439_ _06329_ _06330_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__and2_1
XFILLER_30_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18158_ _08963_ _08997_ _08998_ net337 VGND VGND VPWR VPWR _09006_ sky130_fd_sc_hd__a31oi_4
XPHY_EDGE_ROW_68_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17109_ _07948_ _07977_ _07976_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__nand3_4
X_18089_ _08936_ _08937_ _08903_ VGND VGND VPWR VPWR _08938_ sky130_fd_sc_hd__nand3_2
Xhold369 term_low\[0\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 p_ll\[0\] VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ _09275_ _09384_ _01328_ _01326_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__o31a_1
XFILLER_132_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20051_ net1013 net1043 VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__nand2_1
XFILLER_112_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_146_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_86_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11120_ net697 net517 VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__nand2_1
XFILLER_107_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20318_ net793 net15 VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__and2_1
XFILLER_122_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11051_ net796 _01994_ _01995_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__nor3_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20249_ _01492_ _01447_ net794 _01494_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__o211a_1
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_95_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14810_ net727 net723 net685 net677 VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__nand4_4
X_15790_ _06505_ _06577_ _06664_ _06667_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_4_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11953_ _02886_ _02888_ _02883_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__a21o_1
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _05639_ _05550_ _05463_ _05640_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__and4_4
X_11884_ _02814_ _02819_ _02820_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__o21a_1
X_10904_ net795 net545 net713 VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__and3_1
X_17460_ net340 _08317_ _08321_ _08323_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__nand4_4
X_14672_ _05570_ _05571_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__nand2_2
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16411_ _07223_ _07280_ _07281_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__nand3_2
X_17391_ _08247_ _08248_ _08251_ VGND VGND VPWR VPWR _08258_ sky130_fd_sc_hd__and3_1
X_10835_ p_hl\[30\] net1375 _01847_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__a21oi_1
X_13623_ _04521_ _04522_ _04518_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__a21o_1
X_16342_ _07074_ _07077_ _07075_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_24_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19130_ _10017_ _10019_ net589 net1148 VGND VGND VPWR VPWR _10021_ sky130_fd_sc_hd__nand4_1
X_10766_ p_hl\[22\] p_lh\[22\] VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__and2_1
X_13554_ net1133 _04463_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16273_ _07138_ _07147_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_117_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12505_ _09493_ _09613_ _03258_ _03432_ _03431_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o221ai_2
X_10697_ _01724_ _01728_ _01730_ _01731_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__a211o_1
X_13485_ _04328_ _04394_ _04393_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__o21a_1
XFILLER_9_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19061_ _09937_ _09938_ _09949_ VGND VGND VPWR VPWR _09952_ sky130_fd_sc_hd__nand3_2
XFILLER_138_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12436_ _03365_ _03366_ _03368_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__nand3_1
X_18012_ _04182_ _06441_ _08861_ VGND VGND VPWR VPWR _08862_ sky130_fd_sc_hd__o21ai_4
X_15224_ _06015_ _06032_ _06031_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__o21ai_1
X_15155_ _05997_ _06050_ _06051_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_130_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12367_ net682 net483 VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__nand2_1
X_14106_ net746 net683 VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__nand2_1
X_12298_ _03224_ _03228_ _03229_ _03219_ _03218_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__o2111ai_1
X_11318_ _02257_ _02258_ _09395_ _09613_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19963_ net797 _01186_ _01187_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__nor3b_1
X_15086_ _05980_ _05981_ _05893_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__a21o_1
X_11249_ net697 net1018 net507 net702 VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__a22oi_4
XFILLER_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18914_ _09220_ _09275_ _09801_ VGND VGND VPWR VPWR _09806_ sky130_fd_sc_hd__o21ai_1
X_19894_ net735 net562 net556 net742 VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__a22oi_4
X_14037_ _04913_ _04916_ _04938_ VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__nand3_1
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18845_ _09626_ _09630_ _05044_ _06402_ VGND VGND VPWR VPWR _09737_ sky130_fd_sc_hd__a211o_1
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_128_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ _06862_ _06863_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__nand2_2
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18776_ _09660_ _09661_ _09155_ _09297_ VGND VGND VPWR VPWR _09666_ sky130_fd_sc_hd__o2bb2ai_1
X_17727_ _08588_ _08589_ VGND VGND VPWR VPWR _08590_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_50_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14939_ net726 net723 net677 net864 VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__and4_1
X_17658_ _08517_ _08518_ _08209_ _08376_ VGND VGND VPWR VPWR _08522_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_36_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16609_ _07468_ _07469_ _07474_ _07475_ VGND VGND VPWR VPWR _07481_ sky130_fd_sc_hd__nand4_1
Xclkbuf_leaf_15_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
X_17589_ _08448_ _08450_ _08373_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__and3_1
XFILLER_51_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19328_ net598 net732 _00500_ _00501_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_21_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19259_ net850 _10064_ VGND VGND VPWR VPWR _10160_ sky130_fd_sc_hd__nand2_2
XFILLER_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20103_ _01337_ _01279_ _01336_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__nand3_2
XFILLER_112_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20034_ _01262_ _01263_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__nand2_2
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20798_ clknet_leaf_10_clk _00438_ VGND VGND VPWR VPWR b_h\[4\] sky130_fd_sc_hd__dfxtp_4
X_10620_ net794 net1243 VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__and2_1
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10551_ net793 net1279 VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10482_ _01634_ _01635_ _01641_ _01642_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__a2bb2o_1
Xrebuffer241 net1037 VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlymetal6s2s_1
X_13270_ net923 net766 net710 net704 VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__and4_1
Xrebuffer230 net1025 VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__buf_6
Xrebuffer274 a_l\[9\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd1_1
X_12221_ _03008_ _03151_ net1016 net518 _03150_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o2111ai_4
Xrebuffer263 _05423_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__buf_2
XFILLER_136_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12152_ _02858_ _02925_ _02927_ _02922_ VGND VGND VPWR VPWR _03087_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_112_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11103_ net992 _02044_ _02034_ _02035_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__o211ai_2
X_16960_ _07656_ _07806_ _07825_ _07826_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__nand4_4
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12083_ _03016_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_9_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15911_ a_l\[0\] _06659_ net502 _06660_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__a31o_1
X_11034_ net328 _01977_ _01978_ _01942_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__o211ai_4
XFILLER_110_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16891_ _07759_ net452 _07748_ _07758_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__o211a_1
X_18630_ _09501_ _09502_ _09497_ VGND VGND VPWR VPWR _09507_ sky130_fd_sc_hd__and3_1
X_15842_ _06654_ _06717_ _06716_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__nand3_4
XFILLER_94_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15773_ net239 _06632_ _06633_ _06509_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__a31oi_2
X_18561_ _09430_ _09431_ _09219_ _09222_ VGND VGND VPWR VPWR _09432_ sky130_fd_sc_hd__o2bb2ai_2
X_12985_ _03823_ _03828_ _03829_ VGND VGND VPWR VPWR _03912_ sky130_fd_sc_hd__a21boi_1
X_11936_ _02866_ _02869_ _02870_ _02723_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_92_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17512_ net550 net504 _08209_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__and3_1
X_18492_ net770 net593 VGND VGND VPWR VPWR _09356_ sky130_fd_sc_hd__nand2_1
X_14724_ _05624_ _05610_ _05623_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__nand3_2
XFILLER_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ net565 net494 VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__nand2_1
XFILLER_60_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11867_ _02801_ _02799_ _02800_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__nand3_2
X_14655_ _05553_ _05554_ _05552_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11798_ net637 net546 VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__nand2_1
X_10818_ _01837_ _01832_ net796 VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__a21oi_1
X_17374_ _08199_ _08200_ net234 _08232_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__a22o_1
XFILLER_60_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ _09220_ _09428_ _04508_ _04510_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__o211ai_1
X_14586_ _05472_ _05474_ _05486_ _05487_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__a22o_1
X_16325_ _07193_ _07198_ _07197_ _07189_ VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__o211ai_4
X_10749_ p_hl\[20\] p_lh\[20\] VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__nor2_1
X_19113_ _09727_ _09859_ _09999_ VGND VGND VPWR VPWR _10003_ sky130_fd_sc_hd__o21a_1
X_13537_ _04439_ _04444_ _04445_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand3_2
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16256_ net966 net505 VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19044_ _09931_ _09932_ _09155_ _09340_ VGND VGND VPWR VPWR _09935_ sky130_fd_sc_hd__o2bb2ai_1
X_13468_ _04258_ _04304_ _04305_ _04309_ _04214_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__a32oi_2
X_15207_ _06022_ _06028_ _06100_ _06102_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16187_ _07022_ _07061_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__nand2_1
XFILLER_127_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12419_ a_h\[3\] net474 _03350_ _03351_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__a22o_1
X_13399_ _04308_ _04309_ _04214_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__a21o_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138_ _06012_ _06014_ _06031_ _06033_ VGND VGND VPWR VPWR _06035_ sky130_fd_sc_hd__o211ai_2
X_19946_ _01059_ _01169_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__nand2_1
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15069_ _05963_ _05964_ _05904_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_52_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19877_ net591 net717 _01090_ _01093_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__a22o_1
X_18828_ _09554_ _09556_ _09717_ _09716_ VGND VGND VPWR VPWR _09721_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18759_ _09275_ _09286_ net922 _09639_ _09643_ VGND VGND VPWR VPWR _09648_ sky130_fd_sc_hd__o311a_1
XFILLER_82_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20721_ clknet_leaf_23_clk _00361_ VGND VGND VPWR VPWR p_lh\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20652_ clknet_leaf_12_clk _00292_ VGND VGND VPWR VPWR p_hh\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20583_ clknet_leaf_16_clk _00223_ VGND VGND VPWR VPWR p_hh_pipe\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20017_ _01243_ _01241_ _01245_ VGND VGND VPWR VPWR _01246_ sky130_fd_sc_hd__o21bai_1
XFILLER_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _03696_ _03697_ _03612_ VGND VGND VPWR VPWR _03700_ sky130_fd_sc_hd__a21bo_1
X_11721_ _02482_ _02485_ _02655_ _02656_ _02484_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__o2111ai_1
X_11652_ _01855_ _02589_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__or2_2
X_14440_ net730 net690 VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nand2_1
XFILLER_30_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10603_ _09690_ net1329 VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__and2_1
XFILLER_80_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14371_ _05271_ _05272_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__nand2_2
X_11583_ net681 net510 VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__nand2_1
X_16110_ net1116 net583 net533 net529 VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__nand4_4
X_13322_ net923 net701 VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__nand2_1
X_10534_ net795 net1177 VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__and2_1
X_17090_ net593 net488 _07954_ _07955_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__a22o_1
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10465_ _01626_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__nor2_1
X_16041_ _06858_ _06888_ _06889_ _06913_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__a31oi_2
XFILLER_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13253_ _04160_ _04166_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__nand3_1
X_10396_ _01554_ _01558_ _01562_ _01568_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__a31oi_1
XFILLER_108_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12204_ _03136_ _03137_ _03126_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__nand3_2
X_13184_ _04104_ _04096_ _04103_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__or3_1
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12135_ _03068_ net268 VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19800_ _00912_ _00918_ _00917_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__o21ai_2
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17992_ _08839_ _08841_ _08837_ VGND VGND VPWR VPWR _08843_ sky130_fd_sc_hd__a21o_1
X_16943_ _07810_ _07812_ VGND VGND VPWR VPWR _07813_ sky130_fd_sc_hd__nand2_2
X_12066_ _02895_ _02900_ _02897_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__a21oi_1
X_19731_ _00937_ _00926_ _00898_ _00936_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__o211ai_4
X_11017_ net681 net538 VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__nand2_2
X_16874_ _07740_ _07741_ _09188_ _09668_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19662_ _05044_ _06761_ _00791_ _00819_ _00825_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__o2111ai_4
X_15825_ _06701_ _06703_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__nand2_1
X_18613_ net780 net577 _09480_ _09484_ VGND VGND VPWR VPWR _09488_ sky130_fd_sc_hd__a22o_1
X_19593_ _00789_ net718 net603 _00788_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__and4_4
XFILLER_37_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_125_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _06628_ _06629_ _06575_ VGND VGND VPWR VPWR _06636_ sky130_fd_sc_hd__nand3_2
X_18544_ net737 _09217_ _09410_ _09411_ VGND VGND VPWR VPWR _09413_ sky130_fd_sc_hd__a211o_1
X_12968_ _03893_ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__nand2_1
XFILLER_52_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11919_ _02851_ _02852_ _02853_ _02781_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__o2bb2ai_1
X_15687_ _06455_ _06499_ _06565_ _06566_ VGND VGND VPWR VPWR _06568_ sky130_fd_sc_hd__a2bb2o_1
X_18475_ _09334_ _09335_ net619 net1148 VGND VGND VPWR VPWR _09337_ sky130_fd_sc_hd__and4_1
X_12899_ net645 net1049 net856 net827 VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__and4_1
X_14707_ _05606_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__nand2_1
X_17426_ _08289_ _08290_ _08291_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__a21o_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14638_ _05414_ _05502_ _05503_ _05517_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__a31o_1
X_17357_ _08205_ _08219_ _08220_ VGND VGND VPWR VPWR _08224_ sky130_fd_sc_hd__nand3b_1
X_16308_ _07181_ _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__nand2_1
X_14569_ _05470_ net699 net720 _05469_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__and4_1
XFILLER_118_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17288_ _08008_ _08154_ _08153_ _08152_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__o211ai_4
XFILLER_9_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload20 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_16
Xclkload53 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__inv_8
Xclkload42 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__clkinv_16
X_16239_ net587 net561 net543 net521 VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__nand4_2
Xclkload31 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_41_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19027_ _09915_ _09913_ _09916_ VGND VGND VPWR VPWR _09918_ sky130_fd_sc_hd__nand3_2
XFILLER_127_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19929_ _01146_ _01147_ _01108_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__a21oi_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_50_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20704_ clknet_leaf_34_clk _00344_ VGND VGND VPWR VPWR p_lh\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20635_ clknet_leaf_19_clk _00275_ VGND VGND VPWR VPWR p_hh\[1\] sky130_fd_sc_hd__dfxtp_1
Xclkload3 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_8
X_20566_ clknet_leaf_7_clk _00206_ VGND VGND VPWR VPWR mid_sum\[29\] sky130_fd_sc_hd__dfxtp_1
X_20497_ clknet_leaf_17_clk _00137_ VGND VGND VPWR VPWR term_mid\[41\] sky130_fd_sc_hd__dfxtp_1
X_10250_ _09690_ net1154 VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__and2_1
XFILLER_105_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10181_ net882 VGND VGND VPWR VPWR _09155_ sky130_fd_sc_hd__inv_16
XFILLER_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13940_ net731 net703 VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__nand2_1
XFILLER_115_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15610_ _06470_ _06471_ _06489_ _06490_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__a22o_1
X_13871_ _04629_ _04639_ _04640_ _04641_ _04627_ VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__a32o_1
XFILLER_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16590_ _07459_ _07460_ net814 net1032 VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__nand4_1
XFILLER_74_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12822_ _09493_ _09646_ _03748_ _03749_ VGND VGND VPWR VPWR _03751_ sky130_fd_sc_hd__o211ai_1
X_15541_ _06406_ _06423_ _06424_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__nand3_1
XFILLER_91_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12753_ _03680_ _03682_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__nand2_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _02641_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__inv_2
X_18260_ _08892_ _08947_ _08949_ _09018_ VGND VGND VPWR VPWR _09107_ sky130_fd_sc_hd__nand4_1
X_15472_ _06361_ _06362_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_120_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _08074_ _08077_ _08073_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__o21ai_2
X_12684_ _09439_ _09679_ VGND VGND VPWR VPWR _03614_ sky130_fd_sc_hd__nor2_1
X_14423_ _05318_ _05320_ _05297_ _05298_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__o211ai_2
XFILLER_30_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11635_ _02475_ _02547_ _02545_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__a21o_1
X_18191_ net1119 _09033_ _09035_ VGND VGND VPWR VPWR _09038_ sky130_fd_sc_hd__nand3_4
XFILLER_24_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17142_ _08004_ _08005_ net159 VGND VGND VPWR VPWR _08011_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_96_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _02504_ _02496_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__nand2_1
Xwire630 net632 VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__buf_6
X_14354_ _05100_ _05105_ _05257_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10517_ net1321 _01660_ _01664_ _01666_ net65 VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__a311oi_1
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17073_ _07898_ _07912_ _07916_ _07939_ VGND VGND VPWR VPWR _07942_ sky130_fd_sc_hd__o211ai_1
Xmax_cap418 _07899_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__clkbuf_1
X_13305_ _04192_ _04197_ _04193_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__a21o_1
XFILLER_7_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14285_ _05183_ _05184_ _05033_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__a21oi_1
X_11497_ _02323_ _02223_ net200 VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__a21oi_1
X_16024_ net613 net505 VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__nand2_2
X_13236_ _04145_ _04149_ _04150_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__nand3_1
XFILLER_7_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10448_ _01603_ _01605_ _01609_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__and3_1
X_10379_ _01524_ _01513_ net796 VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__a21oi_1
XFILLER_69_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13167_ _04033_ _04037_ _04067_ _04088_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__o31ai_1
X_12118_ _02836_ _03051_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__nand2_1
X_17975_ net632 net774 _08825_ _08826_ VGND VGND VPWR VPWR _08827_ sky130_fd_sc_hd__a22oi_1
X_13098_ _04019_ _04022_ _04021_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12049_ _02980_ _02974_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__nand2_1
X_16926_ _07792_ _07782_ _07634_ _07794_ VGND VGND VPWR VPWR _07796_ sky130_fd_sc_hd__o211ai_1
X_19714_ _09297_ _00916_ _00919_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__o21ai_2
XFILLER_78_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16857_ _07724_ _07725_ _07727_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__a21o_1
XFILLER_93_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19645_ _00584_ _00587_ _00844_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__o21ai_1
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15808_ _09242_ _09581_ _06440_ _06681_ _06680_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__o221ai_2
X_16788_ net378 _07654_ _07636_ net344 VGND VGND VPWR VPWR _07659_ sky130_fd_sc_hd__o211a_1
XFILLER_80_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19576_ _00766_ _00768_ _00737_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__nand3_2
XFILLER_37_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15739_ net382 _06615_ _06596_ _06614_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_105_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18527_ _09386_ _09393_ VGND VGND VPWR VPWR _09394_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18458_ _09109_ _09208_ _09318_ VGND VGND VPWR VPWR _09320_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_16_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_138_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17409_ _08025_ _08275_ VGND VGND VPWR VPWR _08276_ sky130_fd_sc_hd__nor2_1
X_18389_ _09238_ _09239_ _09234_ VGND VGND VPWR VPWR _09244_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_60_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20420_ clknet_leaf_18_clk _00060_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfxtp_1
X_20351_ net794 net48 VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__and2_1
XFILLER_146_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20282_ net551 net716 VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__nand2_1
XFILLER_130_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11420_ net652 net546 net539 net658 VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__a22oi_1
X_20618_ clknet_leaf_42_clk _00258_ VGND VGND VPWR VPWR p_ll_pipe\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11351_ net678 net519 VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10302_ _00687_ _00698_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__nand2_1
X_20549_ clknet_leaf_54_clk _00189_ VGND VGND VPWR VPWR mid_sum\[12\] sky130_fd_sc_hd__dfxtp_1
X_11282_ _02222_ _02223_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__nor2_1
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070_ net771 net767 net662 net656 VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__and4_1
XFILLER_105_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13021_ _03945_ _03946_ _03878_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__a21o_1
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10233_ net794 net55 VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__and2_1
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17760_ _08278_ _08616_ _08618_ _08273_ VGND VGND VPWR VPWR _08623_ sky130_fd_sc_hd__nand4_2
X_14972_ _05791_ _05868_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__nand2_2
X_16711_ _07433_ _07434_ VGND VGND VPWR VPWR _07582_ sky130_fd_sc_hd__nand2_1
X_17691_ net571 net566 net485 net479 VGND VGND VPWR VPWR _08554_ sky130_fd_sc_hd__and4_1
XFILLER_75_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13923_ _04579_ _04691_ _04581_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_122_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16642_ net939 net948 net523 net570 VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__a22oi_4
XFILLER_90_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13854_ _04752_ _04754_ _04756_ _04740_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__o211ai_4
XFILLER_19_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19430_ net603 net598 net729 net725 VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__nand4_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16573_ _02589_ _06441_ _07317_ _07341_ _07345_ VGND VGND VPWR VPWR _07445_ sky130_fd_sc_hd__o2111ai_2
X_12805_ _03731_ _03733_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__or2_1
X_19361_ _10109_ _10111_ _10070_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__o21ai_2
X_10997_ _01915_ _01923_ _01924_ _01927_ _01914_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__a32oi_4
X_15524_ _09526_ _09581_ _06402_ _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__o31a_1
X_18312_ _09065_ _09146_ _09158_ _09159_ VGND VGND VPWR VPWR _09160_ sky130_fd_sc_hd__o211a_1
X_13785_ _04690_ _04689_ _04688_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__nand3_2
XFILLER_43_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12736_ _03660_ _03662_ _03663_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__a21o_1
X_19292_ _00460_ _00458_ _00461_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _03593_ _03501_ _03592_ _03500_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__a31oi_1
X_18243_ _09040_ _09043_ _09082_ _09083_ VGND VGND VPWR VPWR _09090_ sky130_fd_sc_hd__a22o_1
X_15455_ _06326_ net240 _06327_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_13_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _02553_ _02554_ _02351_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_100_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ _09020_ _09021_ VGND VGND VPWR VPWR _09022_ sky130_fd_sc_hd__nand2_1
X_15386_ _06221_ _06222_ _06225_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__o21ai_1
X_14406_ _09264_ _09460_ _09482_ _05304_ _05303_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__o221a_1
X_17125_ _07947_ _07990_ VGND VGND VPWR VPWR _07994_ sky130_fd_sc_hd__nand2_1
X_12598_ _03513_ _03516_ _03419_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14337_ _05119_ net194 VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__nand2_1
XFILLER_143_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold507 mid_sum\[19\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap226 _03107_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
X_11549_ _02484_ _02486_ net679 net518 VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__nand4_2
Xhold518 mid_sum\[1\] VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap204 _00537_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_1
Xmax_cap259 _07037_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold529 p_lh\[0\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ net561 net509 VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__nand2_2
X_14268_ _05153_ _05154_ _05171_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__o21ai_2
X_16007_ _06537_ _06880_ _06876_ _06879_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__o211a_4
XPHY_EDGE_ROW_115_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13219_ net787 net784 net710 net704 VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__and4_1
X_14199_ _05099_ _05100_ _05103_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__a21bo_1
XFILLER_111_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17958_ net790 net627 net632 net781 VGND VGND VPWR VPWR _08812_ sky130_fd_sc_hd__a22oi_1
X_16909_ _07631_ _07663_ _07778_ VGND VGND VPWR VPWR _07779_ sky130_fd_sc_hd__o21ai_2
X_17889_ _08708_ _08716_ _08746_ VGND VGND VPWR VPWR _08749_ sky130_fd_sc_hd__a21oi_1
X_19628_ _00818_ _00825_ _00823_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_124_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19559_ _00749_ _00742_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__nand2_1
XFILLER_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20403_ clknet_leaf_43_clk _00043_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20334_ net793 net29 VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__and2_2
XPHY_EDGE_ROW_133_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap782 net786 VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__buf_12
X_20265_ _01506_ _01507_ _01508_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_1_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap760 b_l\[6\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__buf_12
Xmax_cap771 net773 VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__buf_12
Xmax_cap793 net795 VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__buf_12
XFILLER_115_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20196_ _01434_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__nor2_1
XFILLER_57_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10920_ net707 net534 VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__nand2_1
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_142_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10851_ net793 net1210 VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__and2_1
XFILLER_72_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10782_ net1349 p_lh\[24\] VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__and2_1
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13570_ _04389_ _04477_ _04479_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__a21o_1
X_12521_ _03158_ _03286_ _03290_ _03450_ VGND VGND VPWR VPWR _03453_ sky130_fd_sc_hd__o211ai_1
XFILLER_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12452_ net674 net489 VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__nand2_1
XFILLER_9_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15240_ _06087_ _06088_ _06130_ _06131_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__a2bb2o_1
X_11403_ _09177_ _09646_ _02339_ _02341_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__o22a_1
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12383_ _03313_ _03315_ _09449_ _09646_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__o2bb2ai_1
X_15171_ _05971_ _05976_ _05979_ _05975_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__a2bb2oi_1
X_11334_ net658 net547 VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__nand2_1
X_14122_ _05019_ _05021_ _05007_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__a21o_1
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11265_ _02199_ net361 net440 VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__nand3_1
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14053_ net157 _04956_ _04958_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__o21bai_4
X_18930_ _09815_ _09817_ _09811_ VGND VGND VPWR VPWR _09822_ sky130_fd_sc_hd__a21o_1
XFILLER_140_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10216_ p_hl\[6\] VGND VGND VPWR VPWR _09537_ sky130_fd_sc_hd__inv_2
X_13004_ _03848_ _03851_ _03807_ _03925_ _03926_ VGND VGND VPWR VPWR _03931_ sky130_fd_sc_hd__a32o_1
X_11196_ _02136_ net180 VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__nor2_1
XFILLER_95_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit202 b_h\[13\] VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__buf_4
X_18861_ _09750_ _09751_ VGND VGND VPWR VPWR _09753_ sky130_fd_sc_hd__nand2_2
XFILLER_121_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit257 a_l\[13\] VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__clkbuf_2
X_17812_ net555 net494 _09373_ VGND VGND VPWR VPWR _08673_ sky130_fd_sc_hd__a21o_1
X_18792_ _09681_ _09682_ VGND VGND VPWR VPWR _09684_ sky130_fd_sc_hd__nand2_1
X_17743_ _08591_ _08592_ _08598_ _08599_ VGND VGND VPWR VPWR _08606_ sky130_fd_sc_hd__nand4_1
X_14955_ _05850_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__nand2_1
X_13906_ _04654_ _04682_ _04806_ _04807_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_18_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17674_ _08533_ _08534_ _08535_ VGND VGND VPWR VPWR _08538_ sky130_fd_sc_hd__a21o_1
X_14886_ _05604_ _05709_ _05712_ _05733_ _05738_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__o2111ai_2
X_19413_ net588 net738 VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__nand2_1
X_16625_ _07355_ _07495_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_102_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13837_ net783 net656 VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__nand2_1
X_16556_ _07421_ _07423_ _07427_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__and3_1
X_13768_ _04669_ net432 _04668_ net286 VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_44_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19344_ _00511_ _00513_ _00519_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__o21ai_1
X_16487_ _07354_ _07356_ a_l\[6\] net502 VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__nand4_2
X_12719_ _03536_ _03540_ _03539_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_15507_ _06394_ _06345_ _06391_ _06393_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__o211ai_1
X_19275_ _10176_ _10164_ _10175_ VGND VGND VPWR VPWR _10177_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_135_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18226_ _08969_ _09059_ _09067_ _09072_ VGND VGND VPWR VPWR _09073_ sky130_fd_sc_hd__o2bb2ai_4
X_15438_ _06326_ _06327_ net241 VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__nand3_1
X_13699_ net762 net683 VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18157_ _08959_ _08960_ _09002_ VGND VGND VPWR VPWR _09005_ sky130_fd_sc_hd__o21ai_1
X_15369_ _06261_ _06262_ net795 VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__o21ai_1
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17108_ net451 _07970_ _07973_ _07964_ _07963_ VGND VGND VPWR VPWR _07977_ sky130_fd_sc_hd__o2111ai_2
X_18088_ _08922_ _08927_ _08929_ _08913_ VGND VGND VPWR VPWR _08937_ sky130_fd_sc_hd__o211ai_2
XFILLER_7_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17039_ _07901_ _07903_ net418 VGND VGND VPWR VPWR _07908_ sky130_fd_sc_hd__a21o_1
XFILLER_89_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold359 p_ll_pipe\[27\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20050_ net568 net1097 VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_146_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20317_ net793 net14 VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap590 a_l\[8\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__buf_8
X_11050_ _01989_ _01991_ _01938_ _01903_ _01940_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__o221a_1
X_20248_ _01491_ _01490_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__nand2_1
XFILLER_131_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20179_ _01415_ _01416_ _01409_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__nand3_2
XFILLER_77_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14740_ _05639_ _05640_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ net653 net647 net526 net520 VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_86_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11883_ _02819_ _02814_ net796 VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_86_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10903_ net794 net1344 VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__and2_1
X_14671_ net750 net655 net649 net756 VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__a22oi_2
X_16410_ net256 _07283_ net257 VGND VGND VPWR VPWR _07284_ sky130_fd_sc_hd__a21oi_2
X_17390_ _08247_ _08248_ _09210_ _09679_ VGND VGND VPWR VPWR _08257_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_83_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10834_ _01849_ _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__or2_1
X_13622_ _09155_ _09460_ _04521_ _04522_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__o211ai_2
X_16341_ _07074_ net484 a_l\[0\] _07075_ VGND VGND VPWR VPWR _07215_ sky130_fd_sc_hd__a31o_1
X_13553_ _04397_ _04459_ _04460_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__nand3_2
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10765_ net795 _01790_ _01791_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__and3_1
X_12504_ _03258_ _03432_ _03428_ _03431_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_43_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19060_ _09938_ _09949_ VGND VGND VPWR VPWR _09951_ sky130_fd_sc_hd__nand2_1
X_16272_ _06962_ _07140_ _07139_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__a21o_1
X_10696_ _01730_ _01731_ _01724_ _01728_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__o211ai_1
X_13484_ net714 net741 _04327_ _04261_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__a22o_1
XFILLER_9_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12435_ _03238_ _03240_ _03239_ VGND VGND VPWR VPWR _03368_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_117_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18011_ _08859_ _08860_ VGND VGND VPWR VPWR _08861_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15223_ _06114_ _06115_ net348 VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__nand3_4
XFILLER_138_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12366_ _03295_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__nand2_1
XFILLER_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15154_ _05998_ _06048_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11317_ _02193_ _02256_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__nand2_2
X_14105_ net746 net683 VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__and2_1
X_12297_ _03224_ _03228_ _03229_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__o21ai_1
X_19962_ _01183_ _01185_ _01182_ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__o21ai_1
X_15085_ _05980_ _05981_ _05893_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__a21oi_1
X_11248_ net698 net510 VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__nand2_1
X_19893_ net742 net735 net563 net556 VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__nand4_2
X_14036_ _04913_ _04916_ _04939_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__a21o_1
X_18913_ _09220_ _09275_ _09801_ VGND VGND VPWR VPWR _09805_ sky130_fd_sc_hd__o21a_1
X_11179_ _02102_ _02119_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__nand2_1
XFILLER_67_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18844_ _09625_ _09629_ _05043_ net847 VGND VGND VPWR VPWR _09736_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_128_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ net1116 net531 net527 a_l\[7\] VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18775_ _09660_ _09661_ net780 net569 VGND VGND VPWR VPWR _09665_ sky130_fd_sc_hd__nand4_2
X_17726_ _08584_ _08586_ _08587_ VGND VGND VPWR VPWR _08589_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_50_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14938_ net723 net677 net866 net726 VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__a22o_1
X_17657_ net416 _08210_ _08518_ _08517_ VGND VGND VPWR VPWR _08521_ sky130_fd_sc_hd__a22oi_1
XFILLER_63_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14869_ _05768_ _05767_ _05766_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__nand3_4
X_16608_ _07468_ _07469_ _07478_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__nand3_1
XFILLER_90_383 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17588_ _08450_ _08373_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__nand2_1
X_19327_ _09231_ _09308_ _00500_ _00501_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__o211ai_1
X_16539_ _07365_ _07366_ _07407_ _07408_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__nand4_2
X_19258_ _10133_ _10119_ _10118_ VGND VGND VPWR VPWR _10159_ sky130_fd_sc_hd__o21ai_2
X_18209_ _09049_ _09055_ VGND VGND VPWR VPWR _09056_ sky130_fd_sc_hd__nor2_1
X_19189_ _10080_ _10082_ VGND VGND VPWR VPWR _10085_ sky130_fd_sc_hd__nand2_1
XFILLER_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20102_ _01280_ _01334_ _01335_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__nand3_2
XFILLER_86_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20033_ _01189_ _01260_ _01261_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__nand3_2
XFILLER_140_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ clknet_leaf_24_clk _00437_ VGND VGND VPWR VPWR b_h\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_10_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ net793 net1293 VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_40_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10481_ _01612_ _01620_ _01628_ _01631_ _01639_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__a41o_1
Xrebuffer220 net1040 VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer231 net1025 VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12220_ _03150_ _03152_ _03148_ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__a21o_1
Xrebuffer242 a_h\[11\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer253 _04513_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__buf_6
Xrebuffer275 a_l\[9\] VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer286 a_l\[4\] VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer297 b_l\[13\] VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd1_1
X_12151_ _02925_ _02858_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_112_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11102_ _02036_ _02045_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__nand2_1
X_12082_ _03009_ _03011_ _03006_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_9_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15910_ _06659_ net502 a_l\[0\] VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__and3_1
X_11033_ net328 _01971_ _01955_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__o21ai_2
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16890_ net452 _07756_ _07747_ _07757_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__o211ai_4
XFILLER_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15841_ _06623_ _06630_ _06714_ _06715_ VGND VGND VPWR VPWR _06720_ sky130_fd_sc_hd__o211ai_2
XFILLER_64_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15772_ _06648_ _06649_ _06650_ net797 VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__a211oi_1
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18560_ _09427_ _09426_ _09324_ VGND VGND VPWR VPWR _09431_ sky130_fd_sc_hd__nand3_4
X_12984_ _03824_ _03825_ _03823_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11935_ _02727_ _02723_ _02726_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o21ai_1
X_17511_ net550 net503 VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__nand2_1
X_18491_ net1124 net585 VGND VGND VPWR VPWR _09355_ sky130_fd_sc_hd__nand2_1
X_14723_ _05618_ net677 net730 VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_28_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _08305_ _08306_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__nand2_1
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14654_ net771 net767 net640 net636 VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__nand4_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11866_ _02802_ _02798_ _02797_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__nand3_4
X_13605_ _04402_ _04507_ _04506_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__o21ai_2
XFILLER_17_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10817_ _01813_ _01833_ _01836_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__a21o_1
X_11797_ net644 net537 VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nand2_1
X_17373_ _08238_ _08237_ _08236_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__nand3_2
X_14585_ net428 _05484_ _05485_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__nand3_2
X_16324_ _07191_ _07192_ _07190_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__o21ai_2
X_10748_ net795 _01775_ _01776_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__and3_1
X_19112_ _09860_ _09998_ _09999_ VGND VGND VPWR VPWR _10002_ sky130_fd_sc_hd__o21ai_2
X_13536_ _04443_ net711 net748 _04442_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__nand4_4
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16255_ net602 net512 net505 net607 VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13467_ _04372_ _04374_ _04266_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__a21o_1
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19043_ _09931_ _09932_ _09929_ VGND VGND VPWR VPWR _09934_ sky130_fd_sc_hd__a21o_1
X_12418_ _03348_ _03210_ _03201_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__nand3b_1
X_10679_ p_hl\[7\] p_lh\[7\] net469 _01715_ VGND VGND VPWR VPWR _01719_ sky130_fd_sc_hd__o211ai_2
X_15206_ _09308_ _09504_ _06097_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__o21ai_1
X_16186_ _07023_ net259 VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__nand2_1
X_13398_ _04214_ _04308_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__nand3_1
Xclone90 net610 VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__clkbuf_16
X_12349_ _03151_ _03279_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__nand2_1
X_15137_ _06026_ _06030_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19945_ _09231_ _09384_ _01060_ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__o21ai_1
X_15068_ _05915_ _05917_ _05960_ _05961_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_52_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net752 net676 VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__nand2_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19876_ _01091_ _01036_ VGND VGND VPWR VPWR _01093_ sky130_fd_sc_hd__nand2_1
XFILLER_95_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18827_ _09716_ _09717_ _09718_ VGND VGND VPWR VPWR _09720_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18758_ _09643_ _09645_ _09639_ VGND VGND VPWR VPWR _09647_ sky130_fd_sc_hd__a21oi_1
X_17709_ _08567_ net490 net1054 _08564_ VGND VGND VPWR VPWR _08572_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_108_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20720_ clknet_leaf_23_clk _00360_ VGND VGND VPWR VPWR p_lh\[22\] sky130_fd_sc_hd__dfxtp_1
X_18689_ _09401_ _09568_ _09563_ _09564_ VGND VGND VPWR VPWR _09572_ sky130_fd_sc_hd__o211ai_4
X_20651_ clknet_leaf_14_clk _00291_ VGND VGND VPWR VPWR p_hh\[17\] sky130_fd_sc_hd__dfxtp_1
X_20582_ clknet_leaf_16_clk _00222_ VGND VGND VPWR VPWR p_hh_pipe\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20016_ _01124_ _01134_ _01121_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__a21o_1
XFILLER_74_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11720_ _02482_ _02485_ _02655_ _02656_ _02484_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_83_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ net486 b_h\[13\] VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__nand2_8
X_10602_ _09690_ net1314 VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__and2_1
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11582_ _02518_ _02481_ _02516_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__nand3_4
X_14370_ net767 net649 net642 net771 VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__a22oi_2
X_10533_ net795 net1181 VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__and2_1
X_13321_ net763 net711 VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nand2_1
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16040_ _06916_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__inv_2
X_10464_ term_mid\[46\] term_high\[46\] VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__nor2_1
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13252_ _04165_ net704 net777 _04164_ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__nand4b_2
X_10395_ term_mid\[35\] term_high\[35\] _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__a21o_1
X_12203_ _09471_ _09613_ _02976_ _03131_ _03130_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__o221ai_4
X_13183_ _04103_ _04104_ _04096_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__o21ai_1
XFILLER_135_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12134_ _03066_ _03060_ _03039_ _03067_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_94_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17991_ _09144_ _09155_ net459 _06521_ _08841_ VGND VGND VPWR VPWR _08842_ sky130_fd_sc_hd__o221ai_1
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19730_ _00937_ _00926_ _00898_ _00936_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__o211a_1
XFILLER_145_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16942_ net554 net550 b_h\[2\] b_h\[3\] VGND VGND VPWR VPWR _07812_ sky130_fd_sc_hd__nand4_4
XFILLER_89_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12065_ _02997_ _02998_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__nand2_1
XFILLER_77_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11016_ _01921_ _01960_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__nand2_4
X_16873_ _02589_ _06605_ net799 net476 _07741_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__o2111ai_4
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19661_ _00787_ _00790_ _00818_ _00824_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__o22ai_2
XFILLER_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15824_ _09188_ _09602_ _06696_ _06697_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__o211ai_1
X_18612_ net780 net576 VGND VGND VPWR VPWR _09487_ sky130_fd_sc_hd__nand2_1
X_19592_ _00785_ _00786_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18543_ _09410_ _09411_ net1082 net737 net847 VGND VGND VPWR VPWR _09412_ sky130_fd_sc_hd__o2111ai_4
X_15755_ _06632_ _06633_ net239 VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__a21oi_2
X_12967_ net976 b_h\[12\] VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__nand2_1
XFILLER_45_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11918_ _02768_ _02782_ _02780_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__a21bo_1
X_15686_ _06565_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__nand2_1
X_18474_ net887 net604 net759 net754 _09330_ VGND VGND VPWR VPWR _09336_ sky130_fd_sc_hd__a41o_1
X_12898_ net645 net638 net856 VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__nand3_2
X_14706_ net720 net1011 _05603_ _05605_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__a22o_1
X_11849_ _02783_ _02768_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__nand2_1
X_17425_ _08052_ _08210_ _08206_ _08208_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14637_ _05509_ _05511_ _05510_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__o21ai_2
X_17356_ _08056_ _08204_ _08219_ _08220_ VGND VGND VPWR VPWR _08223_ sky130_fd_sc_hd__o211ai_2
X_14568_ _05333_ _05467_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__nand2_1
X_16307_ _07050_ _07048_ _07176_ _07178_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__o22ai_4
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17287_ _08006_ _08002_ _08001_ _08014_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__a31oi_1
Xclkload10 clknet_leaf_1_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_2
X_13519_ _04424_ _04426_ _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__o21ai_1
X_14499_ _05110_ _05265_ _05394_ _05399_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__o211ai_1
XFILLER_127_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload43 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__bufinv_16
Xclkload32 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinvlp_4
X_16238_ net561 net522 VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__nand2_2
Xclkload21 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_11_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19026_ net446 _09805_ net368 _09914_ VGND VGND VPWR VPWR _09917_ sky130_fd_sc_hd__o22ai_4
Xclkload54 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__inv_8
X_16169_ _06952_ _07041_ _07042_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__and3_1
XFILLER_127_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19928_ _01030_ _01033_ _01142_ _01143_ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__nand4_1
XFILLER_96_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19859_ _01068_ _01071_ _01073_ VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__nand3_2
XFILLER_52_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ clknet_leaf_34_clk _00343_ VGND VGND VPWR VPWR p_lh\[5\] sky130_fd_sc_hd__dfxtp_1
X_20634_ clknet_leaf_29_clk _00274_ VGND VGND VPWR VPWR p_hh\[0\] sky130_fd_sc_hd__dfxtp_1
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__bufinv_16
XFILLER_137_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20565_ clknet_leaf_7_clk _00205_ VGND VGND VPWR VPWR mid_sum\[28\] sky130_fd_sc_hd__dfxtp_1
X_20496_ clknet_leaf_17_clk _00136_ VGND VGND VPWR VPWR term_mid\[40\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ net622 VGND VGND VPWR VPWR _09144_ sky130_fd_sc_hd__inv_6
XFILLER_59_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13870_ _04629_ _04639_ _04640_ _04641_ _04627_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__a32oi_4
X_12821_ _03748_ _03749_ _03744_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__a21o_1
XFILLER_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15540_ _06421_ _06422_ _06411_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__a21o_1
X_12752_ _03679_ _03522_ _03527_ VGND VGND VPWR VPWR _03682_ sky130_fd_sc_hd__nand3b_1
XFILLER_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _02627_ _02633_ _02632_ net325 _02624_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o2111ai_4
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12683_ _03504_ _03570_ _03573_ _03576_ _03587_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__a32oi_2
XFILLER_70_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15471_ _06358_ net192 _06360_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__or3_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11634_ _02475_ _02547_ _02545_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_120_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _08067_ _08070_ _08076_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__o21ai_1
X_14422_ _05181_ _05321_ _05323_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__nand3_2
XFILLER_15_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18190_ _09030_ _09033_ _09034_ _08987_ VGND VGND VPWR VPWR _09037_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_11_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17141_ _08001_ _08002_ _08006_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _02501_ _02503_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__nand2_1
X_14353_ _05255_ _05256_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__nand2b_1
X_10516_ _01660_ _01664_ net1321 VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__a21oi_1
X_11496_ _02323_ _02223_ net200 VGND VGND VPWR VPWR _02436_ sky130_fd_sc_hd__a21o_1
X_17072_ _07898_ _07912_ _07939_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__o21ai_1
X_13304_ _04200_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__nand2_1
X_14284_ _05177_ _05178_ _05143_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__a21o_1
Xmax_cap408 _00665_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_1
X_10447_ term_mid\[44\] term_high\[44\] VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__xor2_2
X_16023_ _06797_ _06898_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__nand2_2
XFILLER_108_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap419 _07887_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_1
X_13235_ _04149_ _04150_ _04145_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10378_ term_mid\[32\] term_high\[32\] _01482_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__a21o_1
X_13166_ _04033_ _04067_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__nor2_1
X_12117_ net679 net499 net492 net682 VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__a22oi_1
X_17974_ _08824_ _08823_ _08822_ VGND VGND VPWR VPWR _08826_ sky130_fd_sc_hd__nand3_1
X_13097_ _04018_ b_h\[15\] net891 _04017_ _04014_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__a41oi_4
XFILLER_34_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12048_ _09460_ _09613_ _02862_ _02978_ _02977_ VGND VGND VPWR VPWR _02983_ sky130_fd_sc_hd__o221ai_4
X_16925_ _07782_ _07792_ _07634_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__o21ai_2
X_19713_ _00914_ _00915_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__nand2_1
X_19644_ _00844_ _00843_ _00717_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__a21bo_1
X_16856_ net237 _07574_ _07569_ _07572_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__o2bb2ai_2
X_15807_ _06440_ _06681_ net595 net541 _06680_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__o2111ai_2
X_16787_ _07656_ _07636_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__nand2_1
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19575_ _00734_ _00736_ net273 _00767_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__o22ai_4
X_13999_ _04746_ _04890_ _04900_ _04902_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__a2bb2oi_2
X_15738_ net1008 _06595_ _06617_ VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_105_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18526_ _09246_ _09352_ _09389_ _09390_ VGND VGND VPWR VPWR _09393_ sky130_fd_sc_hd__o211ai_2
X_18457_ _09098_ net149 _09317_ _09104_ VGND VGND VPWR VPWR _09318_ sky130_fd_sc_hd__o22ai_2
XFILLER_61_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17408_ _08020_ _08021_ _08156_ _08158_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__nand4_1
X_15669_ net309 _06533_ _06546_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_16_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18388_ _09233_ net371 _09241_ VGND VGND VPWR VPWR _09243_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_60_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17339_ net566 net503 VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20350_ net794 net47 VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__and2_1
X_19009_ _09872_ _09898_ _09899_ VGND VGND VPWR VPWR _09900_ sky130_fd_sc_hd__nand3_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20281_ _01502_ _01525_ _01527_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__a21oi_1
XFILLER_114_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20617_ clknet_leaf_42_clk _00257_ VGND VGND VPWR VPWR p_ll_pipe\[15\] sky130_fd_sc_hd__dfxtp_1
X_11350_ net1078 net517 VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_78_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20548_ clknet_leaf_42_clk _00188_ VGND VGND VPWR VPWR mid_sum\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10301_ term_low\[22\] term_mid\[22\] VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__nand2_1
X_11281_ _02115_ _02117_ _02220_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__a21oi_4
X_13020_ _03878_ _03946_ VGND VGND VPWR VPWR _03947_ sky130_fd_sc_hd__nand2_1
X_20479_ clknet_leaf_45_clk _00119_ VGND VGND VPWR VPWR term_mid\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10232_ net794 net44 VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_109_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16710_ _07434_ _07441_ _07581_ _07579_ net797 VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__a311oi_1
XFILLER_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14971_ _05789_ _05790_ _05867_ _05868_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__a22o_1
X_17690_ net566 net479 VGND VGND VPWR VPWR _08553_ sky130_fd_sc_hd__nand2_1
X_13922_ _04826_ _04821_ _04825_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__a21o_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16641_ net939 net947 VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_89_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13853_ _04736_ _04737_ _04752_ _04754_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__o22ai_2
X_16572_ _07315_ _07316_ _07341_ _07345_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12804_ _03728_ _03729_ _03730_ _03673_ VGND VGND VPWR VPWR _03733_ sky130_fd_sc_hd__o211a_1
X_19360_ _00488_ _00490_ _00528_ _00529_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__nand4_2
X_10996_ _01927_ _01914_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__nand2_1
X_15523_ _06406_ _06407_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__nand2_1
X_18311_ _09150_ _09151_ _09155_ _09242_ VGND VGND VPWR VPWR _09159_ sky130_fd_sc_hd__o2bb2ai_1
X_13784_ _04689_ _04688_ _04690_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__a21o_1
XFILLER_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12735_ _03660_ _03662_ _03663_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__a21oi_1
XFILLER_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19291_ _00458_ _00460_ net1148 net579 VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__nand4_2
X_12666_ _03596_ _03500_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__nand2_1
X_18242_ _09082_ _09083_ net277 VGND VGND VPWR VPWR _09089_ sky130_fd_sc_hd__a21oi_1
X_15454_ _06217_ _06340_ _06344_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_13_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _02448_ _02548_ _02549_ _02352_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__a31oi_2
XTAP_TAPCELL_ROW_100_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _08943_ _08945_ _09016_ _09017_ VGND VGND VPWR VPWR _09021_ sky130_fd_sc_hd__o211ai_2
X_12597_ _03525_ _03419_ _03522_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__nand3_2
X_15385_ _09504_ _09515_ net455 _06225_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__o31a_1
X_14405_ _05303_ _05306_ _05301_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__a21o_1
X_11548_ _09449_ _09602_ _02483_ _02485_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__o22ai_2
X_17124_ _07947_ _07986_ _07987_ _07989_ VGND VGND VPWR VPWR _07993_ sky130_fd_sc_hd__a31oi_2
X_14336_ _05186_ _05190_ _05228_ _05230_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__o2bb2ai_2
Xhold508 p_hh\[26\] VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xwire483 b_h\[12\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__buf_8
Xmax_cap205 _10130_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xmax_cap238 _06853_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_133_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11479_ _02389_ _02390_ _02416_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17055_ _07784_ _07923_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__nand2_2
Xhold519 term_mid\[16\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ _05168_ _05170_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__nand2_2
X_16006_ _06879_ _06882_ _06876_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__a21oi_4
XFILLER_124_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13218_ _01855_ net459 _04135_ net795 VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__o211a_1
X_14198_ _04694_ _04829_ _04964_ net142 _05101_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__o41a_1
X_13149_ a_h\[13\] _04043_ b_h\[14\] _04041_ _04047_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a311oi_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17957_ _09690_ net632 net790 VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__and3_1
X_16908_ _07664_ _07690_ VGND VGND VPWR VPWR _07778_ sky130_fd_sc_hd__nand2_2
X_17888_ _08715_ _08712_ _08709_ _08747_ VGND VGND VPWR VPWR _08748_ sky130_fd_sc_hd__a211oi_1
XFILLER_66_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclone351 b_l\[8\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__clkbuf_16
X_16839_ net629 net472 _07707_ _07709_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__a22oi_2
XFILLER_53_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19627_ _00817_ _00819_ _00822_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__nand3_2
XFILLER_81_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19558_ _00746_ _00748_ _00743_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__a21oi_1
X_18509_ net791 net782 net577 net569 VGND VGND VPWR VPWR _09375_ sky130_fd_sc_hd__nand4_2
XFILLER_21_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19489_ _00643_ _00645_ _00667_ _00669_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__nand4_4
XFILLER_147_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20402_ clknet_leaf_43_clk _00042_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfxtp_1
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20333_ net795 net28 VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__and2_1
XFILLER_103_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap772 net773 VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__buf_12
X_20264_ net724 net551 b_l\[14\] net548 VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__nand4_1
Xmax_cap761 net762 VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__buf_12
Xmax_cap794 _09690_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_73_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap783 net786 VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__buf_8
X_20195_ _01429_ _01432_ _01425_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10850_ net793 net1211 VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__and2_1
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10781_ net795 _01804_ _01805_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__and3_1
X_12520_ _03425_ net322 _03447_ VGND VGND VPWR VPWR _03452_ sky130_fd_sc_hd__nand3b_2
XFILLER_52_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ net674 net489 VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__and2_1
XFILLER_138_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11402_ net712 net487 VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__nand2_1
X_15170_ _06058_ _06060_ _06063_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__nand3_1
X_12382_ net672 net665 net995 net492 VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__nand4_2
XFILLER_4_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14121_ _05019_ _05021_ _05007_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__a21oi_1
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11333_ net671 net536 VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__nand2_1
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11264_ _02199_ net361 net440 VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_115_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14052_ _04811_ _04815_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__nand2_1
X_10215_ net547 VGND VGND VPWR VPWR _09526_ sky130_fd_sc_hd__inv_4
XFILLER_97_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13003_ _03848_ _03851_ _03807_ _03925_ _03926_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__a32oi_2
X_18860_ net603 net1091 net737 net609 VGND VGND VPWR VPWR _09752_ sky130_fd_sc_hd__a22oi_1
X_11195_ _02055_ _01991_ _02056_ net213 VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__o31ai_4
X_17811_ _08632_ _08633_ _08638_ _08639_ VGND VGND VPWR VPWR _08672_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18791_ net760 net596 net1001 net1111 VGND VGND VPWR VPWR _09683_ sky130_fd_sc_hd__a22oi_2
Xsplit236 b_l\[10\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__buf_2
X_17742_ _08592_ _08598_ _08599_ VGND VGND VPWR VPWR _08605_ sky130_fd_sc_hd__nand3_1
XFILLER_0_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14954_ _05691_ _05847_ _05851_ net311 VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__o211ai_4
X_17673_ _08533_ _08534_ _08535_ VGND VGND VPWR VPWR _08537_ sky130_fd_sc_hd__nand3_1
X_13905_ _04811_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__inv_2
X_16624_ net1069 net513 net506 net590 VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__a22oi_4
X_14885_ _05604_ _05709_ _05712_ _05733_ _05738_ VGND VGND VPWR VPWR _05784_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_18_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19412_ net591 net732 VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__nand2_2
X_13836_ net778 net660 VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__nand2_2
X_16555_ _07421_ _07423_ _07427_ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__a21oi_2
X_10979_ _09406_ _09592_ _01887_ _01921_ _01920_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_102_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13767_ _04671_ _04670_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_44_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19343_ _00519_ _00516_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__nand2_1
X_16486_ _09231_ _09613_ _07357_ _07358_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__o211ai_2
X_12718_ _03536_ _03539_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__nand2_1
XFILLER_71_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15506_ _06341_ _06343_ _06394_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__a21oi_1
X_19274_ _09220_ _09319_ _10172_ VGND VGND VPWR VPWR _10176_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_135_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18225_ _09061_ _09066_ VGND VGND VPWR VPWR _09072_ sky130_fd_sc_hd__nand2_2
X_15437_ _06326_ _06327_ net241 VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__a21o_1
X_13698_ _04520_ _04589_ _04600_ _04601_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_135_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ net682 net679 net483 net481 _03402_ VGND VGND VPWR VPWR _03580_ sky130_fd_sc_hd__a41o_1
XFILLER_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18156_ _09000_ _09001_ _08961_ VGND VGND VPWR VPWR _09004_ sky130_fd_sc_hd__nand3_1
X_15368_ _06208_ _06216_ _06217_ _06210_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__a31oi_1
X_17107_ _07963_ _07964_ _07971_ _07972_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__o2bb2ai_1
X_18087_ _08910_ net374 _08930_ VGND VGND VPWR VPWR _08936_ sky130_fd_sc_hd__o21ai_2
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14319_ _05024_ _05221_ _05222_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nand3_4
X_15299_ _02362_ net455 _06119_ _06123_ _06193_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__o2111ai_2
X_17038_ _07906_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18989_ _09749_ _09754_ _09752_ VGND VGND VPWR VPWR _09880_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_146_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone170 net687 VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__clkbuf_16
XFILLER_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20316_ net793 net13 VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__and2_1
Xmax_cap580 net581 VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__buf_12
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20247_ _01487_ _01489_ _01451_ _01455_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__o22ai_1
Xmax_cap591 net592 VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__buf_8
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20178_ _01415_ _01416_ _09373_ _01408_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_76_326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11951_ net1016 net524 VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11882_ _02815_ _02816_ _02569_ _02691_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10902_ net794 net1348 VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__and2_1
X_14670_ net750 net655 VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__nand2_1
X_10833_ p_hl\[31\] p_lh\[31\] VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__and2_1
X_13621_ _04524_ _04525_ _04527_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__nand3_2
X_16340_ _07206_ _07207_ _07211_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__nand3_2
X_10764_ _01778_ _01787_ _01789_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__o21ai_1
X_13552_ _04457_ _04458_ _04398_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12503_ _09493_ _09613_ _03434_ VGND VGND VPWR VPWR _03435_ sky130_fd_sc_hd__o21ai_1
X_16271_ _07145_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__inv_2
X_18010_ net623 net774 VGND VGND VPWR VPWR _08860_ sky130_fd_sc_hd__nand2_1
X_10695_ p_hl\[11\] p_lh\[11\] VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__nand2_1
X_13483_ _04329_ _04330_ _04392_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__a21o_1
XFILLER_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12434_ _03239_ _03243_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15222_ net348 _06116_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__nand3b_4
X_12365_ _03294_ _03296_ _03297_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__nand3_4
X_15153_ _05916_ _05962_ _06046_ _06047_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_130_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11316_ net698 net691 net1018 net507 VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__nand4_2
X_19961_ _01179_ _01181_ _01183_ _01185_ VGND VGND VPWR VPWR _01186_ sky130_fd_sc_hd__a211oi_1
XFILLER_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15084_ _05893_ _05980_ _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__nand3_1
X_14104_ _04874_ _04877_ _04878_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__a21o_1
XFILLER_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12296_ _03224_ _03228_ _03229_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__o21a_1
X_14035_ _04936_ net317 _04909_ _04915_ _04913_ VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__o221ai_4
X_18912_ net446 _09800_ _09798_ VGND VGND VPWR VPWR _09804_ sky130_fd_sc_hd__o21bai_1
XFILLER_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11247_ net708 net501 VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__nand2_1
XFILLER_4_396 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19892_ net742 net735 net563 VGND VGND VPWR VPWR _01111_ sky130_fd_sc_hd__nand3_1
X_11178_ _02095_ _02100_ _02119_ _02099_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__o211ai_2
XFILLER_94_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18843_ _09731_ _09732_ _09735_ net794 VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__o211a_1
XFILLER_67_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18774_ _09155_ _09297_ _09660_ _09661_ VGND VGND VPWR VPWR _09664_ sky130_fd_sc_hd__o211ai_1
X_15986_ net1116 net531 VGND VGND VPWR VPWR _06863_ sky130_fd_sc_hd__nand2_1
X_17725_ _08577_ _08585_ _08580_ _08583_ _08587_ VGND VGND VPWR VPWR _08588_ sky130_fd_sc_hd__o221ai_4
XFILLER_48_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14937_ net723 net677 net861 net726 VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__a22oi_4
XFILLER_36_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17656_ _08210_ _08518_ net416 _08517_ VGND VGND VPWR VPWR _08520_ sky130_fd_sc_hd__nand4_4
X_14868_ _05549_ _05644_ _05643_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__o21a_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16607_ _07468_ _07469_ _07476_ _07477_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o2bb2ai_1
X_17587_ _08448_ _08450_ _08373_ VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__a21o_1
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13819_ _04719_ _04721_ _04722_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__and3_1
XFILLER_23_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16538_ _07407_ _07408_ _07367_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__a21o_1
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14799_ _05692_ _05693_ _05695_ net807 VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__o2bb2ai_1
X_19326_ _00500_ _00501_ _00496_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__a21o_1
X_16469_ _07338_ _07340_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__nand3_1
X_19257_ _10140_ _10143_ _10141_ VGND VGND VPWR VPWR _10157_ sky130_fd_sc_hd__a21boi_4
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18208_ net774 net610 net769 net605 _09048_ VGND VGND VPWR VPWR _09055_ sky130_fd_sc_hd__a41o_1
X_19188_ _10079_ _10081_ VGND VGND VPWR VPWR _10084_ sky130_fd_sc_hd__nor2_1
XFILLER_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18139_ net774 net971 net769 net615 VGND VGND VPWR VPWR _08987_ sky130_fd_sc_hd__a22oi_1
XFILLER_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20101_ _01324_ _01329_ _01330_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__nand3_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20032_ _01188_ _01159_ _01258_ _01259_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__o211ai_4
XFILLER_112_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20796_ clknet_leaf_24_clk _00436_ VGND VGND VPWR VPWR b_h\[2\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_81_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_40_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10480_ _01595_ _01616_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__a21o_1
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer210 _06596_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__buf_1
Xrebuffer232 _01252_ VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer254 _06592_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__buf_6
Xrebuffer243 a_h\[11\] VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd1_1
X_12150_ _03035_ _03037_ _03081_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__nand3_2
Xrebuffer276 _01262_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__buf_1
Xrebuffer298 b_l\[13\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__buf_8
X_11101_ _02042_ _02044_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_112_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12081_ _09493_ _09602_ _02884_ _03007_ _03011_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_9_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11032_ _01954_ _01972_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__nand2_1
XFILLER_77_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15840_ _06623_ _06630_ _06716_ _06717_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_1_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15771_ _06501_ _06568_ _06647_ _06460_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__and4_1
XFILLER_85_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12983_ _03908_ net885 net645 _03906_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__nand4_4
X_11934_ _02628_ _02722_ _02727_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__o21a_1
X_17510_ _09373_ _09613_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__nor2_1
XFILLER_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18490_ net764 net597 VGND VGND VPWR VPWR _09354_ sky130_fd_sc_hd__nand2_1
X_14722_ _09308_ _09449_ _05479_ _05616_ _05615_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__o221ai_2
XFILLER_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17441_ net565 net498 net493 net569 VGND VGND VPWR VPWR _08307_ sky130_fd_sc_hd__a22oi_2
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14653_ net771 net767 net640 net636 VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_28_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _02669_ _02604_ _02672_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__o21a_1
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13604_ _04510_ _04508_ _04506_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__a21o_1
X_10816_ p_hl\[27\] p_lh\[27\] _01834_ _01835_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__a211o_1
X_11796_ net646 net535 VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__nand2_1
X_17372_ _08079_ _08082_ _08136_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__o21ai_1
X_19111_ _09865_ _10000_ _10001_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__o21a_1
X_14584_ net428 _05482_ _05483_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__nand3b_2
X_16323_ _07194_ _07196_ _07190_ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__a21o_1
X_10747_ _01766_ _01772_ _01774_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__o21ai_1
X_13535_ _04440_ net701 net757 VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__nand3_1
XFILLER_139_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16254_ net602 net513 VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10678_ _01710_ _01715_ net469 VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__a21oi_1
X_13466_ _04264_ _04263_ _04374_ _04372_ VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__o211ai_1
X_19042_ _09155_ _09340_ _09931_ _09932_ VGND VGND VPWR VPWR _09933_ sky130_fd_sc_hd__o211ai_2
X_12417_ _03202_ _03348_ _03349_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__nand3_1
X_15205_ _06094_ _06096_ _06098_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__a21oi_2
X_16185_ _06845_ _07058_ _07053_ _07057_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__o2bb2ai_4
X_13397_ _04306_ _04307_ _04257_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__nand3_2
XFILLER_142_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12348_ net633 net526 net1023 net1036 VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__a22oi_2
X_15136_ _06024_ _06025_ _06016_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nand3_1
X_12279_ _03206_ _03208_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__nand2_1
X_19944_ _01160_ _01162_ _01086_ VGND VGND VPWR VPWR _01168_ sky130_fd_sc_hd__nand3_2
X_15067_ _05959_ _05956_ _05918_ _05916_ _05958_ VGND VGND VPWR VPWR _05965_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_52_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14018_ net752 net683 net676 net758 VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__a22o_1
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19875_ _01037_ _01089_ _01088_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__a21oi_1
X_18826_ _09716_ _09717_ _09718_ VGND VGND VPWR VPWR _09719_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_143_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15969_ _06748_ _06823_ _06821_ net261 VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_110_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18757_ net775 net770 net581 net576 VGND VGND VPWR VPWR _09645_ sky130_fd_sc_hd__nand4_1
XFILLER_82_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17708_ _08566_ _08570_ VGND VGND VPWR VPWR _08571_ sky130_fd_sc_hd__nor2_1
X_18688_ _09326_ _09397_ _09398_ _09403_ _09422_ VGND VGND VPWR VPWR _09571_ sky130_fd_sc_hd__a32oi_1
XTAP_TAPCELL_ROW_108_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17639_ _08396_ _08402_ _08498_ _08499_ VGND VGND VPWR VPWR _08503_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_23_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20650_ clknet_leaf_14_clk _00290_ VGND VGND VPWR VPWR p_hh\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20581_ clknet_leaf_16_clk _00221_ VGND VGND VPWR VPWR p_hh_pipe\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_63_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19309_ _10179_ _10162_ _00475_ _00473_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__o211ai_2
XFILLER_32_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20015_ _01099_ _01239_ _01103_ _01237_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__nand4_4
XFILLER_48_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11650_ net486 b_h\[13\] VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__and2_4
XFILLER_23_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20779_ clknet_leaf_22_clk _00419_ VGND VGND VPWR VPWR a_l\[1\] sky130_fd_sc_hd__dfxtp_4
X_11581_ _02481_ _02516_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__nand2_1
X_10601_ net794 net1200 VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__and2_1
X_10532_ net795 net1175 VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__and2_1
XFILLER_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13320_ _04231_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__nand2_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10463_ term_mid\[46\] term_high\[46\] VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__and2_1
X_13251_ _04163_ _04165_ _04161_ VGND VGND VPWR VPWR _04166_ sky130_fd_sc_hd__o21ai_1
X_10394_ term_mid\[35\] term_high\[35\] term_mid\[34\] term_high\[34\] VGND VGND VPWR
+ VPWR _01567_ sky130_fd_sc_hd__o211a_1
X_12202_ _03130_ _03132_ _03133_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__a21o_1
X_13182_ _04078_ _04100_ _04101_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__and3_1
X_12133_ _03038_ _03064_ _03065_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_94_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17990_ net781 net615 net611 net790 VGND VGND VPWR VPWR _08841_ sky130_fd_sc_hd__a22o_1
XFILLER_89_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12064_ _02997_ _02998_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__and2_1
X_16941_ net550 net530 VGND VGND VPWR VPWR _07811_ sky130_fd_sc_hd__nand2_1
XFILLER_145_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11015_ net681 net947 VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__nand2_1
XFILLER_104_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16872_ _07741_ net476 net798 _07740_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__and4_1
XFILLER_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19660_ _00787_ _00790_ _00818_ _00824_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__o22a_1
X_15823_ _06692_ _06696_ _06697_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__and3_1
XFILLER_65_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18611_ _09155_ _09286_ VGND VGND VPWR VPWR _09486_ sky130_fd_sc_hd__nor2_1
X_19591_ net598 net591 net729 net725 VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__nand4_2
XFILLER_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _06631_ _06623_ net239 _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__o211ai_4
XFILLER_80_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18542_ _09166_ _09308_ _04555_ _06441_ _09408_ VGND VGND VPWR VPWR _09411_ sky130_fd_sc_hd__o221a_1
X_12966_ net873 net999 VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__nand2_1
XFILLER_46_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14705_ _05467_ _05604_ net720 net1011 _05603_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__o2111ai_4
X_11917_ _02766_ _02767_ _02780_ VGND VGND VPWR VPWR _02853_ sky130_fd_sc_hd__o21a_1
X_15685_ _06496_ _06558_ _06559_ _06561_ VGND VGND VPWR VPWR _06566_ sky130_fd_sc_hd__nand4_2
X_18473_ net609 net604 net759 net754 VGND VGND VPWR VPWR _09335_ sky130_fd_sc_hd__nand4_1
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12897_ net638 net856 VGND VGND VPWR VPWR _03825_ sky130_fd_sc_hd__nand2_1
X_11848_ _02766_ _02767_ _02780_ _02782_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__a2bb2o_1
X_17424_ _08288_ net503 net1004 _08287_ VGND VGND VPWR VPWR _08290_ sky130_fd_sc_hd__nand4_4
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14636_ _05412_ _05521_ _05522_ _05524_ _05526_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__a32oi_2
X_17355_ _08054_ _08062_ _08219_ _08220_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__a22o_1
XFILLER_60_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14567_ net727 net723 net695 net690 VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__nand4_1
XFILLER_14_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16306_ _07051_ _07177_ _07179_ VGND VGND VPWR VPWR _07181_ sky130_fd_sc_hd__nand3b_4
X_11779_ _02713_ _02702_ _02712_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__nand3_1
X_13518_ _04411_ _04421_ _04422_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__nand3_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17286_ _08004_ _08005_ net159 _08013_ VGND VGND VPWR VPWR _08154_ sky130_fd_sc_hd__a31oi_2
X_14498_ _05110_ _05265_ _05394_ _05399_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__o211a_1
X_19025_ _09798_ net446 _09801_ VGND VGND VPWR VPWR _09916_ sky130_fd_sc_hd__o21ai_1
X_16237_ net561 net543 net521 net587 VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__a22o_1
Xclkload44 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinv_8
Xclkload33 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinv_4
Xclkload11 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__inv_6
XFILLER_62_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13449_ _04353_ _04357_ _04358_ _04345_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__o211ai_1
Xclkload22 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_11_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__inv_6
X_16168_ _07038_ _07040_ _06951_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_11_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15119_ _05925_ _05929_ _05928_ VGND VGND VPWR VPWR _06016_ sky130_fd_sc_hd__o21ai_1
X_16099_ _06875_ _06887_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__nand2_1
XFILLER_87_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19927_ _01142_ _01144_ VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__nand2_1
X_19858_ _01072_ _01074_ VGND VGND VPWR VPWR _01075_ sky130_fd_sc_hd__nand2_1
X_18809_ net1031 net1081 _09695_ _09696_ VGND VGND VPWR VPWR _09702_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19789_ _00996_ _00998_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__nor2_1
XFILLER_70_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20702_ clknet_leaf_39_clk _00342_ VGND VGND VPWR VPWR p_lh\[4\] sky130_fd_sc_hd__dfxtp_1
X_20633_ clknet_leaf_49_clk _00273_ VGND VGND VPWR VPWR p_ll_pipe\[31\] sky130_fd_sc_hd__dfxtp_1
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__bufinv_16
XFILLER_20_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20564_ clknet_leaf_17_clk _00204_ VGND VGND VPWR VPWR mid_sum\[27\] sky130_fd_sc_hd__dfxtp_1
X_20495_ clknet_leaf_27_clk _00135_ VGND VGND VPWR VPWR term_mid\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12820_ net648 net645 b_h\[9\] net828 VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__nand4_2
XFILLER_28_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12751_ _03680_ VGND VGND VPWR VPWR _03681_ sky130_fd_sc_hd__inv_2
X_11702_ _02625_ _02637_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__nand2_1
X_12682_ _03583_ _03584_ _03582_ VGND VGND VPWR VPWR _03612_ sky130_fd_sc_hd__a21bo_1
X_15470_ _06358_ net192 _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__o21ai_1
X_11633_ _02439_ _02560_ _02562_ _02569_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_120_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14421_ net931 _05321_ _05323_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__nand3_4
X_17140_ _08006_ _08002_ _08001_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_96_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ net652 net646 net546 net537 VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__nand4_4
Xwire610 net611 VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__buf_12
X_14352_ _05253_ _05096_ _05254_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__nand3_2
XFILLER_10_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10515_ net793 _01663_ _01665_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__and3_1
X_11495_ _02433_ _02434_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__nand2_1
X_17071_ _07914_ _07915_ _07936_ _07938_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__o22ai_2
X_13303_ _04189_ _04201_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__nand2_1
X_14283_ _05139_ _05141_ _05178_ _05177_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__o211ai_2
Xmax_cap409 _00600_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_1
X_10446_ _01609_ _01610_ _01611_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__o21a_1
X_16022_ net613 net512 net505 net1127 VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__a22oi_2
Xwire687 net688 VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__buf_12
X_13234_ _01871_ _04134_ net777 net710 _04148_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__o2111ai_1
XFILLER_6_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10377_ term_mid\[33\] term_high\[33\] VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__xor2_2
XFILLER_124_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13165_ _04031_ _04065_ _04066_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__o21ai_1
XFILLER_124_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12116_ net679 net499 VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__nand2_1
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17973_ _08822_ _08823_ _08824_ VGND VGND VPWR VPWR _08825_ sky130_fd_sc_hd__a21o_1
X_13096_ _04012_ _04013_ _04019_ _04020_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a22oi_1
XFILLER_2_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12047_ _02862_ _02978_ net1048 net501 _02977_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__o2111ai_2
X_16924_ _07783_ _07786_ _07780_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__a21o_1
X_19712_ net574 net1033 net567 net834 VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__a22oi_4
X_16855_ _07725_ VGND VGND VPWR VPWR _07726_ sky130_fd_sc_hd__inv_2
X_19643_ _00840_ _00841_ _00720_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__nand3_2
X_15806_ _06680_ _06683_ _09242_ _09581_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16786_ net378 _07654_ net344 VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__o21ai_1
X_19574_ _00766_ _00768_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__nand2_1
XFILLER_34_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13998_ _04748_ _04889_ _04900_ _04902_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__o211ai_4
X_15737_ net382 _06615_ _06614_ VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_105_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12949_ _03875_ _03876_ net793 VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o21ai_1
X_18525_ _09246_ _09352_ _09383_ _09385_ VGND VGND VPWR VPWR _09392_ sky130_fd_sc_hd__a2bb2oi_1
X_15668_ net309 _06533_ _06546_ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__a21oi_1
X_18456_ _09202_ _09204_ _09019_ VGND VGND VPWR VPWR _09317_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_47_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17407_ _08023_ _08160_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__nor2_2
XFILLER_61_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14619_ _05513_ _05515_ _05506_ _05507_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_16_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15599_ net625 net616 net531 net527 VGND VGND VPWR VPWR _06481_ sky130_fd_sc_hd__nand4_4
X_18387_ net459 _07100_ net780 net585 _09238_ VGND VGND VPWR VPWR _09241_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_60_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17338_ net571 _08054_ net503 _08056_ VGND VGND VPWR VPWR _08205_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_60_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17269_ _08084_ _08086_ _08128_ _08130_ VGND VGND VPWR VPWR _08137_ sky130_fd_sc_hd__nand4_1
X_19008_ _09895_ _09879_ VGND VGND VPWR VPWR _09899_ sky130_fd_sc_hd__nand2_1
X_20280_ _01525_ _01502_ net794 VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20616_ clknet_leaf_42_clk _00256_ VGND VGND VPWR VPWR p_ll_pipe\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20547_ clknet_leaf_42_clk _00187_ VGND VGND VPWR VPWR mid_sum\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11280_ _02115_ _02117_ _02220_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__and3_1
XFILLER_125_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10300_ term_low\[22\] term_mid\[22\] VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__or2_1
XFILLER_106_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10231_ net794 net33 VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__and2_1
X_20478_ clknet_leaf_45_clk _00118_ VGND VGND VPWR VPWR term_mid\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_109_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14970_ _05789_ _05790_ _05867_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_109_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13921_ _04826_ _04821_ _04825_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__a21oi_2
XFILLER_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16640_ net572 net516 VGND VGND VPWR VPWR _07512_ sky130_fd_sc_hd__nand2_1
X_13852_ _04758_ _04740_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__nand2_2
X_16571_ _07420_ _07422_ _07421_ _07426_ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__a22oi_2
X_12803_ _03673_ _03730_ _03729_ _03728_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__a211o_1
X_13783_ _04688_ _04689_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__a21oi_1
X_10995_ _01938_ _01903_ net795 _01940_ _01939_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__o2111a_1
X_15522_ net625 net1105 _06404_ _06405_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__a22o_1
X_12734_ _03549_ _03555_ _03556_ _03547_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__a31o_1
X_18310_ _09150_ _09151_ net779 net593 VGND VGND VPWR VPWR _09158_ sky130_fd_sc_hd__nand4_1
XFILLER_55_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19290_ _00458_ _00460_ b_l\[8\] net579 VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_54_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_8
X_18241_ _09082_ _09083_ _09044_ VGND VGND VPWR VPWR _09088_ sky130_fd_sc_hd__nand3_1
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12665_ _03588_ _03595_ _03594_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__o21ai_1
X_15453_ _06301_ _06305_ _06335_ _06342_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_13_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11616_ _02553_ _02554_ _02348_ _02350_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_100_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18172_ _09015_ net218 _09014_ VGND VGND VPWR VPWR _09020_ sky130_fd_sc_hd__nand3_4
X_12596_ _03521_ _03517_ _03420_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__a21oi_1
X_14404_ _05303_ _05306_ _05301_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__a21oi_1
X_15384_ _06275_ _06276_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__nand2_1
Xwire440 _02202_ VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_1
X_17123_ _07990_ _07991_ VGND VGND VPWR VPWR _07992_ sky130_fd_sc_hd__nand2_1
X_11547_ net671 net664 net525 net520 VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__nand4_2
X_14335_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__inv_2
XFILLER_116_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold509 p_lh\[26\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
X_17054_ net561 net514 VGND VGND VPWR VPWR _07923_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_133_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16005_ net602 net572 net543 net521 VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__nand4_2
X_11478_ _02389_ _02390_ _02416_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__nand3_1
XFILLER_109_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14266_ _05165_ _05160_ net429 net391 VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__o211ai_4
X_10429_ term_mid\[41\] term_high\[41\] VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__nor2_1
X_13217_ net784 net713 net707 net1088 VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__a22o_1
X_14197_ _04828_ _04962_ _04963_ _04695_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nand4_4
X_13148_ _04054_ b_h\[15\] net869 _04052_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__a31o_1
XFILLER_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17956_ _08810_ _08811_ net796 VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13079_ net641 net1149 net1112 a_h\[13\] VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_29_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone330 net620 VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__clkbuf_16
X_16907_ _07775_ _07776_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__nand2_2
X_17887_ _08746_ VGND VGND VPWR VPWR _08747_ sky130_fd_sc_hd__inv_2
X_16838_ _07473_ _07474_ _07483_ _07487_ VGND VGND VPWR VPWR _07709_ sky130_fd_sc_hd__nand4_1
X_19626_ _00817_ _00822_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__nand2_2
X_16769_ net936 net903 VGND VGND VPWR VPWR _07640_ sky130_fd_sc_hd__nand2_4
X_19557_ _00748_ net567 b_l\[8\] _00746_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__nand4_2
X_18508_ _09370_ _09371_ VGND VGND VPWR VPWR _09374_ sky130_fd_sc_hd__nand2_1
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_22_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19488_ _00643_ _00645_ _00666_ _00668_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_34_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18439_ _09223_ _09224_ _09290_ _09295_ _09296_ VGND VGND VPWR VPWR _09299_ sky130_fd_sc_hd__o221ai_4
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_38_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20401_ clknet_leaf_46_clk _00041_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfxtp_1
XFILLER_147_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20332_ net793 net27 VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__and2_1
XFILLER_107_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap762 net763 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__buf_8
Xmax_cap773 net775 VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__buf_12
Xmax_cap751 net752 VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__buf_6
X_20263_ net551 b_l\[14\] net548 net724 VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__a22o_1
XFILLER_143_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap784 net785 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__buf_12
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20194_ _01433_ _01434_ _01425_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__o21ba_1
XFILLER_142_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_47_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_96_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_37_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10780_ _01792_ _01799_ _01803_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__o21ai_1
XFILLER_12_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12450_ _03309_ _03315_ net460 VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11401_ net706 net975 net492 net708 VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__a22oi_2
XFILLER_40_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12381_ net665 net495 VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__nand2_1
X_14120_ _05008_ _05019_ _05021_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__and3_1
X_11332_ net362 _02177_ _02176_ VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__a21boi_2
XFILLER_141_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11263_ _02199_ net440 VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_115_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14051_ _04799_ _04800_ _04952_ _04953_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__o211ai_4
X_11194_ _02129_ _02130_ _02135_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__nand3_2
XFILLER_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13002_ _03807_ _03852_ _03925_ _03926_ VGND VGND VPWR VPWR _03929_ sky130_fd_sc_hd__nand4_1
X_10214_ net907 VGND VGND VPWR VPWR _09515_ sky130_fd_sc_hd__inv_6
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17810_ _08669_ net130 _08671_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__o21a_1
XFILLER_95_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18790_ net760 net596 VGND VGND VPWR VPWR _09682_ sky130_fd_sc_hd__nand2_1
XFILLER_94_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17741_ _08593_ _08600_ _08601_ VGND VGND VPWR VPWR _08604_ sky130_fd_sc_hd__nand3_1
X_14953_ _05833_ _05834_ _05842_ _05843_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__o2bb2ai_1
X_17672_ _08535_ VGND VGND VPWR VPWR _08536_ sky130_fd_sc_hd__inv_2
XFILLER_48_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13904_ _04810_ _04702_ _04809_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__nand3_2
X_14884_ _05749_ _05760_ _05761_ _05750_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__a31o_1
X_16623_ net584 net513 VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__nand2_2
XFILLER_90_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13835_ _04592_ _04595_ _04597_ VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_18_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19411_ _00496_ _00501_ _00499_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__a21oi_2
XFILLER_35_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_90_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16554_ _07213_ _07425_ _07424_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__o21bai_1
X_10978_ _01887_ _01921_ net697 net1106 _01920_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_102_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13766_ _04499_ _04501_ _04670_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_44_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19342_ _00518_ _00505_ _00507_ _00517_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__o211ai_1
X_16485_ _07262_ net513 net590 VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__nand3_1
X_12717_ _09482_ _09646_ _03639_ _09635_ _03642_ VGND VGND VPWR VPWR _03647_ sky130_fd_sc_hd__o221ai_2
X_15505_ _06365_ _06384_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__or2_1
X_13697_ _04591_ _04598_ _04520_ _04589_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__o2bb2ai_4
X_19273_ _10168_ _10171_ net765 net562 VGND VGND VPWR VPWR _10175_ sky130_fd_sc_hd__nand4_2
X_12648_ _03576_ _03578_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__nand2_1
X_18224_ _09066_ _09068_ _09061_ VGND VGND VPWR VPWR _09071_ sky130_fd_sc_hd__a21oi_2
X_15436_ _09384_ _09493_ _06280_ _06282_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_135_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18155_ _09000_ _09001_ _08961_ VGND VGND VPWR VPWR _09003_ sky130_fd_sc_hd__and3_1
X_17106_ net451 _07970_ _07973_ VGND VGND VPWR VPWR _07975_ sky130_fd_sc_hd__o21a_1
X_12579_ _03506_ _03508_ b_h\[8\] VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__nand3_1
X_15367_ _06258_ _06260_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__nand2_1
XFILLER_117_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18086_ _08880_ _08865_ _08879_ _08931_ _08932_ VGND VGND VPWR VPWR _08935_ sky130_fd_sc_hd__o2111ai_4
X_15298_ _06009_ _06107_ _09362_ _09471_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__a211o_1
X_14318_ _05216_ _05198_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__nand2_1
X_17037_ _07899_ _07901_ _07903_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__nand3_2
X_14249_ net761 net662 _05151_ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_55_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18988_ _09873_ _09876_ _09878_ VGND VGND VPWR VPWR _09879_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17939_ _09373_ _09679_ _08782_ VGND VGND VPWR VPWR _08796_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_146_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19609_ net409 _00794_ _00803_ _00804_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__o211ai_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_18_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20315_ net793 net11 VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__and2_1
Xmax_cap570 net571 VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__buf_8
Xmax_cap581 net584 VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_55_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20246_ _01443_ _01446_ _01451_ _01455_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__o22ai_1
Xmax_cap592 net596 VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__buf_12
XFILLER_107_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20177_ _01369_ _01410_ net1013 net721 _01414_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__o2111ai_4
XFILLER_130_273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11950_ _02725_ _02884_ VGND VGND VPWR VPWR _02886_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ net794 net1335 VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__and2_1
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11881_ _02565_ _02567_ _02691_ _02441_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_86_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10832_ p_hl\[31\] p_lh\[31\] VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__nor2_1
XFILLER_60_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13620_ _04524_ _04525_ _04527_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__and3_1
X_10763_ p_hl\[20\] p_lh\[20\] _01779_ _01785_ _01789_ VGND VGND VPWR VPWR _01790_
+ sky130_fd_sc_hd__a221o_1
X_13551_ _04458_ _04457_ _04398_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nand3_4
XFILLER_53_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16270_ _07138_ net345 _07141_ VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__o21ai_2
X_12502_ _03261_ _03430_ _03432_ _03258_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10694_ p_hl\[11\] p_lh\[11\] VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__and2_1
X_13482_ net714 net741 VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nand2_2
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15221_ _06103_ _06106_ _06113_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12433_ _03224_ _03227_ _03357_ _03360_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_117_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12364_ _03273_ _03275_ _03289_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_73_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15152_ _05916_ _05962_ _06046_ _06047_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__and4_2
XFILLER_141_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11315_ net691 net510 VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__nand2_1
XFILLER_99_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19960_ _00975_ _00976_ _01184_ VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15083_ _05977_ _05978_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__nand2_1
X_14103_ _04707_ _04923_ _04926_ _04922_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_130_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12295_ _03223_ _03224_ _03226_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14034_ _04936_ net317 _04909_ _04915_ _04913_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__o221a_1
X_18911_ net446 _09801_ net763 net580 VGND VGND VPWR VPWR _09803_ sky130_fd_sc_hd__nand4b_1
X_11246_ _02063_ _02068_ _02065_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__a21oi_1
X_19891_ net742 net556 VGND VGND VPWR VPWR _01110_ sky130_fd_sc_hd__nand2_2
X_11177_ _02099_ _02101_ _02119_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__a21o_1
XFILLER_122_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18842_ _09437_ _09584_ _09728_ _09734_ VGND VGND VPWR VPWR _09735_ sky130_fd_sc_hd__o31a_1
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15985_ a_l\[7\] net527 VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__nand2_1
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18773_ _09662_ _09655_ VGND VGND VPWR VPWR _09663_ sky130_fd_sc_hd__nand2_1
XFILLER_94_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17724_ _08488_ _08503_ _08502_ VGND VGND VPWR VPWR _08587_ sky130_fd_sc_hd__o21ai_2
X_14936_ net720 net685 VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_128_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17655_ _08513_ _08516_ _08479_ VGND VGND VPWR VPWR _08519_ sky130_fd_sc_hd__a21boi_1
X_14867_ _05748_ _05750_ _05763_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_141_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16606_ _07474_ _07475_ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__nand2_1
X_17586_ _08448_ _08450_ _08373_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13818_ _04722_ _04721_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__nand2_1
X_14798_ _05692_ _05693_ _05694_ _05572_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16537_ net1030 _07367_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__nand2_1
X_13749_ _04656_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__inv_2
XFILLER_16_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19325_ net591 net588 net744 net738 VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__nand4_4
X_16468_ _07335_ _07312_ _07334_ VGND VGND VPWR VPWR _07341_ sky130_fd_sc_hd__nand3_2
X_19256_ _10007_ _10138_ _10139_ _10141_ _10144_ VGND VGND VPWR VPWR _10156_ sky130_fd_sc_hd__a32oi_2
XTAP_TAPCELL_ROW_42_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16399_ _07258_ _07270_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__and3_1
X_18207_ _09049_ _09051_ _09048_ VGND VGND VPWR VPWR _09054_ sky130_fd_sc_hd__o21ai_1
X_19187_ net621 net718 _10077_ _10078_ VGND VGND VPWR VPWR _10082_ sky130_fd_sc_hd__a22o_1
X_15419_ net726 net722 net640 net635 VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__nand4_1
XFILLER_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18138_ net615 net774 net971 net769 VGND VGND VPWR VPWR _08986_ sky130_fd_sc_hd__nand4_4
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18069_ net781 net605 VGND VGND VPWR VPWR _08918_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_7_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
X_20100_ _01331_ _01323_ _01321_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_70_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20031_ _01198_ _01194_ _01197_ _01254_ _01256_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__o2111ai_2
XFILLER_85_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20795_ clknet_leaf_23_clk _00435_ VGND VGND VPWR VPWR b_h\[1\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_81_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer211 _06593_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__buf_1
Xrebuffer200 _02510_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_20_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer233 _07408_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__buf_2
XFILLER_108_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer299 net1095 VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer277 _00645_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer288 b_l\[1\] VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__buf_1
XFILLER_135_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11100_ _01948_ _01944_ _02039_ _02038_ _01947_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__o221a_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12080_ _02884_ _03007_ net906 net518 _03011_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_9_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11031_ net328 _01971_ _01954_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20229_ _01422_ _01470_ _01418_ _01419_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__nand4_2
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15770_ _06645_ _06646_ _06649_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__a21oi_2
X_12982_ _03906_ _03908_ _09515_ _09646_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11933_ _09449_ _09613_ _02867_ _02868_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o211ai_2
XFILLER_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14721_ _05611_ _05619_ _05620_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__nand3_1
XFILLER_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11864_ _02604_ net952 _02672_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__o21ai_1
X_17440_ net565 net498 VGND VGND VPWR VPWR _08306_ sky130_fd_sc_hd__nand2_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14652_ net767 net640 net636 net771 VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_28_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ p_hl\[27\] p_lh\[27\] p_hl\[26\] p_lh\[26\] VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__o211a_1
X_17371_ _08135_ _08130_ _08083_ VGND VGND VPWR VPWR _08238_ sky130_fd_sc_hd__a21oi_1
XFILLER_72_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13603_ _04510_ net689 net762 _04508_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__and4_1
X_16322_ net620 net812 net496 net491 VGND VGND VPWR VPWR _07196_ sky130_fd_sc_hd__nand4_1
X_11795_ _02612_ _02616_ VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__nand2_1
X_19110_ _09865_ _10000_ net797 VGND VGND VPWR VPWR _10001_ sky130_fd_sc_hd__a21oi_1
X_14583_ _05480_ _05481_ net730 net685 VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__nand4_1
XFILLER_13_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10746_ _01766_ _01772_ _01774_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__or3_1
X_13534_ _04441_ net705 net751 VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__nand3_1
X_16253_ _06993_ _07012_ _07121_ _07122_ VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__o211ai_4
X_10677_ p_hl\[8\] p_lh\[8\] VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__xor2_1
X_13465_ _04372_ _04374_ _04265_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nand3_1
X_19041_ b_l\[0\] net1086 net552 net549 VGND VGND VPWR VPWR _09932_ sky130_fd_sc_hd__nand4_4
XFILLER_145_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16184_ _07058_ _06845_ _07053_ _07057_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__o2bb2a_1
X_12416_ _03201_ _03203_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__nand2_1
X_15204_ _06094_ _06096_ _06098_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__nand3_2
X_13396_ _04258_ _04304_ _04305_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__nand3_1
X_15135_ _06024_ _06025_ _06016_ VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__and3_1
XFILLER_142_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12347_ net637 net633 net526 net524 VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__nand4_2
XFILLER_142_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12278_ _03209_ _03211_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__nand2_1
X_19943_ _01166_ VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__inv_2
X_15066_ _05956_ _05959_ _05915_ _05917_ _05958_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__o221ai_1
X_11229_ net671 net664 net547 net539 VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__nand4_2
XFILLER_68_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19874_ _01037_ _01039_ _01088_ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14017_ net758 net676 VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__nand2_1
X_18825_ _09547_ _09550_ _09551_ _09556_ VGND VGND VPWR VPWR _09718_ sky130_fd_sc_hd__a31o_1
XFILLER_83_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15968_ _06733_ _06836_ _06738_ _06842_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__o22ai_4
XFILLER_83_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18756_ net775 net1146 net580 net576 VGND VGND VPWR VPWR _09644_ sky130_fd_sc_hd__and4_1
X_15899_ _06774_ _06775_ net613 net515 VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__and4_1
X_17707_ _08564_ net490 a_l\[13\] VGND VGND VPWR VPWR _08570_ sky130_fd_sc_hd__nand3_1
X_18687_ _09403_ _09422_ VGND VGND VPWR VPWR _09569_ sky130_fd_sc_hd__nand2_1
XFILLER_48_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14919_ _05815_ _05814_ _05811_ _05816_ VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__o22ai_1
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17638_ _08398_ _08489_ _08498_ _08499_ VGND VGND VPWR VPWR _08502_ sky130_fd_sc_hd__o211ai_2
XFILLER_63_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17569_ net585 net581 _02588_ _08320_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__a31o_1
X_20580_ clknet_leaf_17_clk _00220_ VGND VGND VPWR VPWR p_hh_pipe\[10\] sky130_fd_sc_hd__dfxtp_1
X_19308_ net298 _00452_ _00472_ _00474_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_63_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19239_ _10128_ net205 _10118_ _10120_ VGND VGND VPWR VPWR _10139_ sky130_fd_sc_hd__o211ai_2
XFILLER_117_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20014_ _01238_ _01105_ _01235_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__nor3_2
XFILLER_101_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10600_ _09690_ net1165 VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__and2_1
X_20778_ clknet_leaf_22_clk _00418_ VGND VGND VPWR VPWR a_l\[0\] sky130_fd_sc_hd__dfxtp_4
X_11580_ _02369_ _02480_ _02515_ _02514_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__o211ai_4
XFILLER_23_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10531_ net795 net1241 VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__and2_1
XFILLER_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13250_ net784 net700 net693 net787 VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__a22oi_2
X_10462_ _01617_ _01620_ _01612_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__a31oi_1
XFILLER_109_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12201_ _02976_ _03131_ net665 net501 _03130_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__o2111ai_4
X_10393_ _01417_ _01513_ _01554_ net470 VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nand4_1
XFILLER_124_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13181_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__inv_2
X_12132_ _03063_ _03047_ VGND VGND VPWR VPWR _03067_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_94_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16940_ _07645_ _07809_ VGND VGND VPWR VPWR _07810_ sky130_fd_sc_hd__nand2_1
X_12063_ net637 net633 net537 net535 VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__nand4_4
X_11014_ net691 net534 VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__nand2_1
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16871_ _07738_ _07739_ VGND VGND VPWR VPWR _07741_ sky130_fd_sc_hd__nand2_1
X_15822_ _06696_ _06697_ _06692_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__a21o_1
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18610_ _09480_ _09484_ VGND VGND VPWR VPWR _09485_ sky130_fd_sc_hd__nand2_1
X_19590_ net598 net591 _05043_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_125_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15753_ _06627_ _06584_ VGND VGND VPWR VPWR _06633_ sky130_fd_sc_hd__nand2_4
X_12965_ net1015 net976 b_h\[12\] b_h\[13\] VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__nand4_1
X_18541_ _09405_ _09408_ _09409_ VGND VGND VPWR VPWR _09410_ sky130_fd_sc_hd__a21oi_2
XFILLER_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11916_ _02826_ _02849_ _02850_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__nand3_2
X_14704_ net727 net723 net690 net685 VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__nand4_1
X_15684_ _06554_ _06556_ _06562_ _06557_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__o211ai_1
XFILLER_73_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18472_ _09331_ _09332_ VGND VGND VPWR VPWR _09334_ sky130_fd_sc_hd__nand2_1
X_12896_ net645 net823 VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__nand2_1
X_11847_ _02768_ _02780_ _02782_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__nand3_1
X_17423_ net1004 net503 _08287_ _08288_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__a22o_1
X_14635_ net65 _05535_ _05536_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__nor3_1
X_11778_ _02710_ _02711_ _02703_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__a21oi_1
X_17354_ _08219_ _08220_ _08205_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__a21oi_2
X_14566_ net727 net723 net695 net689 VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__and4_1
XFILLER_14_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16305_ _07050_ _07177_ _07179_ _07047_ VGND VGND VPWR VPWR _07180_ sky130_fd_sc_hd__and4b_1
X_17285_ _08140_ _08146_ _08149_ _08145_ VGND VGND VPWR VPWR _08153_ sky130_fd_sc_hd__o211ai_4
X_10729_ net468 _01756_ _01758_ net796 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a31o_1
X_13517_ _04423_ _04425_ _04410_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__nand3_1
XFILLER_14_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16236_ net561 net1063 net521 net590 VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__a22oi_4
X_14497_ _05110_ _05265_ _05394_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__o21ai_1
X_19024_ net457 _06985_ net592 net748 _09910_ VGND VGND VPWR VPWR _09915_ sky130_fd_sc_hd__o2111ai_1
Xclkload34 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload34/X sky130_fd_sc_hd__clkbuf_8
Xclkload23 clknet_leaf_40_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_16
X_13448_ _04353_ _04357_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__o21ai_1
Xclkload12 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_11_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16167_ _07041_ _07042_ _06952_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__a21oi_1
Xclkload45 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__inv_12
X_13379_ _09155_ _09428_ _04222_ _04287_ _04286_ VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__o221ai_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16098_ _06972_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__nand2_2
X_15118_ _06012_ _06014_ VGND VGND VPWR VPWR _06015_ sky130_fd_sc_hd__nor2_1
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19926_ _01142_ _01143_ net295 VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__a21o_1
X_15049_ _05944_ a_h\[7\] net719 _05943_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__and4_1
XFILLER_130_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19857_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__inv_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18808_ _09688_ _09692_ _09694_ VGND VGND VPWR VPWR _09701_ sky130_fd_sc_hd__nand3_1
X_19788_ _00888_ _00889_ net407 _00995_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__a31o_1
XFILLER_83_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18739_ _09595_ _09621_ _09623_ VGND VGND VPWR VPWR _09626_ sky130_fd_sc_hd__nand3_4
XFILLER_49_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20701_ clknet_leaf_39_clk _00341_ VGND VGND VPWR VPWR p_lh\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20632_ clknet_leaf_49_clk _00272_ VGND VGND VPWR VPWR p_ll_pipe\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20563_ clknet_leaf_17_clk _00203_ VGND VGND VPWR VPWR mid_sum\[26\] sky130_fd_sc_hd__dfxtp_1
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_4
XFILLER_109_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20494_ clknet_leaf_18_clk _00134_ VGND VGND VPWR VPWR term_mid\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12750_ _03528_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__nand2_1
XFILLER_43_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11701_ _02627_ _02636_ _02635_ net325 _02624_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__o2111ai_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12681_ _03502_ _03589_ _03591_ _03594_ _03500_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__a32o_1
X_11632_ _02566_ _02568_ _02570_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_120_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _05316_ _05317_ _05297_ _05298_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__o211ai_2
X_14351_ _05253_ _05254_ _05096_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a21oi_1
XFILLER_128_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ net872 net855 VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__nand2_4
X_13302_ _04213_ _04214_ VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__nand2_1
X_10514_ _01653_ _01657_ _01664_ term_high\[55\] VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__nand4_2
X_11494_ _02247_ _02430_ _02432_ VGND VGND VPWR VPWR _02434_ sky130_fd_sc_hd__nand3b_2
X_17070_ _07785_ _07919_ _07934_ net343 VGND VGND VPWR VPWR _07939_ sky130_fd_sc_hd__o211ai_2
XFILLER_7_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire655 net657 VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__buf_6
X_14282_ _05033_ _05184_ _05183_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__nand3_4
X_10445_ _01610_ _01609_ net796 VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__a21oi_1
X_16021_ net613 net512 VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__nand2_2
XFILLER_109_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13233_ net777 net710 _04147_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__a22o_1
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13164_ _04070_ _04085_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__xnor2_2
X_10376_ _01417_ _01460_ _01493_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__o21a_1
X_12115_ net687 net489 VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__nand2_1
XFILLER_2_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17972_ _09155_ _09166_ _08814_ _06441_ net459 VGND VGND VPWR VPWR _08824_ sky130_fd_sc_hd__o32ai_2
X_13095_ _04018_ b_h\[15\] net838 _04017_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nand4_1
X_12046_ _09460_ _09613_ _02980_ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__o21ai_1
X_16923_ _07783_ _07786_ _07780_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__a21oi_1
X_19711_ net1079 net574 net1033 net567 VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__nand4_1
X_16854_ _07718_ _07720_ _07722_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__nand3_1
X_19642_ _00721_ _00837_ _00839_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__nand3_2
XFILLER_38_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15805_ _06680_ _06683_ _09242_ _09581_ VGND VGND VPWR VPWR _06684_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16785_ _07653_ _07643_ _07638_ _07651_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__o211ai_4
XFILLER_92_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19573_ net367 _00756_ _00760_ net406 VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__o211ai_2
X_13997_ _04748_ _04889_ _04900_ _04902_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__o211a_1
X_15736_ _06524_ _06527_ _06610_ _06611_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__nand4_1
X_12948_ _03786_ _03794_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__nand2_1
X_18524_ _09246_ _09352_ _09390_ VGND VGND VPWR VPWR _09391_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15667_ net309 _06533_ net346 VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_105_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18455_ net153 _09312_ _09315_ VGND VGND VPWR VPWR _09316_ sky130_fd_sc_hd__a21o_1
X_12879_ _03507_ b_h\[8\] net633 VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_47_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17406_ _08156_ _08272_ VGND VGND VPWR VPWR _08273_ sky130_fd_sc_hd__nand2_2
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14618_ _05506_ _05507_ _05513_ _05515_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_16_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15598_ net1100 net803 VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__nand2_8
X_18386_ _09238_ _09239_ _09155_ _09253_ VGND VGND VPWR VPWR _09240_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_138_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17337_ _08054_ net503 net571 VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14549_ _09220_ _09504_ _05447_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__o21ai_1
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17268_ _08086_ _08128_ _08130_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__nand3_2
X_16219_ net570 net541 VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__and2_1
X_17199_ _08060_ _08065_ _08063_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__o21a_1
X_19007_ _09877_ _09878_ _09890_ _09894_ VGND VGND VPWR VPWR _09898_ sky130_fd_sc_hd__o211ai_2
XFILLER_6_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19909_ net589 net721 _01126_ _01129_ VGND VGND VPWR VPWR _01130_ sky130_fd_sc_hd__a22oi_2
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20615_ clknet_leaf_41_clk _00255_ VGND VGND VPWR VPWR p_ll_pipe\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20546_ clknet_leaf_43_clk _00186_ VGND VGND VPWR VPWR mid_sum\[9\] sky130_fd_sc_hd__dfxtp_1
X_10230_ net797 VGND VGND VPWR VPWR _09690_ sky130_fd_sc_hd__clkinv_16
X_20477_ clknet_leaf_47_clk _00117_ VGND VGND VPWR VPWR term_mid\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_91_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13920_ _04693_ _04824_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nor2_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13851_ _04752_ _04754_ _04756_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__o21ai_2
X_16570_ _07420_ _07422_ _07421_ _07426_ VGND VGND VPWR VPWR _07442_ sky130_fd_sc_hd__a22o_1
X_10994_ _01901_ _01938_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__or2_1
X_12802_ _03673_ _03730_ _03729_ _03728_ VGND VGND VPWR VPWR _03731_ sky130_fd_sc_hd__a211oi_1
X_13782_ _04393_ _04570_ _04573_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__o21ai_2
XFILLER_43_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15521_ _06404_ _06405_ net625 net1105 VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__nand4_2
X_12733_ _03549_ _03555_ _03556_ _03547_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__a31oi_2
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18240_ _08999_ _09006_ _09085_ _09086_ VGND VGND VPWR VPWR _09087_ sky130_fd_sc_hd__o211ai_4
X_15452_ _06301_ _06305_ _06335_ _06342_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__o31a_1
X_12664_ _03502_ _03591_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__nand2_1
X_14403_ net756 net750 net667 net662 VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_13_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _02448_ _02548_ _02549_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_100_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18171_ _09015_ net218 _09014_ VGND VGND VPWR VPWR _09019_ sky130_fd_sc_hd__and3_1
X_12595_ net353 _03517_ _03519_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__nand3_1
X_15383_ _06271_ _06272_ _06273_ _06233_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__a22o_1
Xwire441 _01856_ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_2
X_11546_ net672 net664 net526 net520 VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__and4_1
X_17122_ _07983_ _07984_ _07987_ _07947_ VGND VGND VPWR VPWR _07991_ sky130_fd_sc_hd__o211ai_4
XFILLER_7_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14334_ _05232_ _05234_ _05186_ _05190_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__o211ai_2
Xwire430 _04882_ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_1
XFILLER_144_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17053_ net578 net503 VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__nand2_1
Xmax_cap207 _09095_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
X_14265_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__inv_2
Xwire496 net497 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_133_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16004_ net966 net572 net1063 net521 VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__and4_1
X_11477_ _02389_ _02390_ _02414_ _02415_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__o2bb2ai_1
Xmax_cap218 net219 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
X_13216_ net792 net786 VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__nand2_8
X_10428_ _01590_ _01595_ _01596_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__o21a_1
X_14196_ _04822_ _04959_ _04961_ _04962_ _04827_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__a32oi_4
X_13147_ _04017_ _04059_ _04060_ _04061_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a31o_1
XFILLER_3_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10359_ _01161_ _01300_ _01289_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__o21a_1
X_17955_ _09373_ _09668_ _08780_ _08796_ _08798_ VGND VGND VPWR VPWR _08811_ sky130_fd_sc_hd__o32a_1
X_13078_ a_h\[13\] net641 net1152 net1112 VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__nand4_1
X_12029_ _02819_ _02814_ _02812_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__a21o_1
X_16906_ _07772_ _07770_ _07766_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__nand3b_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17886_ _08743_ _08745_ VGND VGND VPWR VPWR _08746_ sky130_fd_sc_hd__nand2_1
Xclone331 net627 VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__clkbuf_16
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16837_ _07473_ _07474_ _07483_ _07487_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__and4_1
XFILLER_81_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19625_ _00783_ _00815_ _00816_ _00821_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__a31oi_2
X_16768_ net936 net904 VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__and2_1
X_19556_ _00746_ _00748_ _09264_ _09297_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_19_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15719_ net602 net541 VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__and2_1
X_18507_ net782 net577 net569 net791 VGND VGND VPWR VPWR _09372_ sky130_fd_sc_hd__a22oi_4
X_16699_ _07564_ _07565_ _07450_ VGND VGND VPWR VPWR _07571_ sky130_fd_sc_hd__a21o_1
X_19487_ _00643_ _00645_ _00671_ _00673_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__nand4_2
X_18438_ _09290_ _09295_ _09296_ VGND VGND VPWR VPWR _09298_ sky130_fd_sc_hd__o21ai_2
XFILLER_22_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18369_ _09221_ VGND VGND VPWR VPWR _09222_ sky130_fd_sc_hd__inv_2
XFILLER_147_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20400_ clknet_leaf_46_clk _00040_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20331_ net793 net26 VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20262_ _09340_ _09384_ _01503_ _01505_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__o22a_1
Xmax_cap741 net742 VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_8
Xmax_cap763 net765 VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__buf_12
Xmax_cap752 net753 VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__buf_12
XFILLER_103_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap774 net1123 VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__clkbuf_8
X_20193_ _01430_ _01431_ _01426_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__a21oi_1
Xmax_cap796 net65 VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__buf_12
Xmax_cap785 net786 VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_102_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ net708 net706 net975 net492 VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__nand4_1
X_12380_ _03310_ _03311_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__nand2_1
XFILLER_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11331_ _02176_ _02179_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__nand2_1
XFILLER_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20529_ clknet_leaf_47_clk _00169_ VGND VGND VPWR VPWR term_low\[24\] sky130_fd_sc_hd__dfxtp_1
X_11262_ _02199_ net361 _02201_ net464 VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_118_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14050_ _04799_ _04800_ _04952_ _04953_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__o211a_1
X_11193_ _02129_ _02130_ _02135_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__and3_1
XFILLER_133_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13001_ _03856_ _03927_ VGND VGND VPWR VPWR _03928_ sky130_fd_sc_hd__nor2_1
X_10213_ net651 VGND VGND VPWR VPWR _09504_ sky130_fd_sc_hd__clkinv_8
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17740_ _08591_ _08592_ _08600_ _08601_ VGND VGND VPWR VPWR _08603_ sky130_fd_sc_hd__nand4_1
XFILLER_0_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14952_ _05840_ _05841_ _05833_ _05834_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__o211ai_2
X_17671_ _08432_ _08437_ _08436_ VGND VGND VPWR VPWR _08535_ sky130_fd_sc_hd__a21bo_1
X_13903_ _04774_ _04776_ _04800_ _04802_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__o2bb2ai_1
X_14883_ _05670_ _05744_ _05745_ _05760_ _05761_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__a32oi_4
X_16622_ net950 net503 VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__nand2_1
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19410_ _00496_ _00501_ _00499_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__a21o_1
X_13834_ _04738_ _04739_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nor2_1
XFILLER_46_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19341_ _00505_ _00518_ _00507_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__o21ai_1
X_16553_ _07213_ _07425_ _07424_ VGND VGND VPWR VPWR _07426_ sky130_fd_sc_hd__o21ba_1
X_10977_ net697 net1106 _01920_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__a22o_2
XFILLER_90_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13765_ net432 _04669_ _04668_ _04671_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_44_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16484_ _07353_ net506 a_l\[7\] VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__nand3_1
X_12716_ _03643_ _03635_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__nand2_1
X_15504_ _06392_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__inv_2
X_13696_ _04603_ _04590_ _04602_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__nand3_4
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19272_ _10172_ net562 net765 VGND VGND VPWR VPWR _10174_ sky130_fd_sc_hd__nand3_1
X_12647_ _03504_ _03570_ _03573_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__nand3_2
X_18223_ net459 _06867_ net779 net1113 _09068_ VGND VGND VPWR VPWR _09070_ sky130_fd_sc_hd__o2111ai_4
X_15435_ _06325_ _06288_ _06324_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_135_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18154_ _09000_ _09001_ VGND VGND VPWR VPWR _09002_ sky130_fd_sc_hd__nand2_1
X_15366_ net150 _06257_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__nand2_1
X_17105_ net451 _07970_ _07973_ VGND VGND VPWR VPWR _07974_ sky130_fd_sc_hd__o21ai_2
X_12578_ _03432_ _03505_ _03507_ _03430_ VGND VGND VPWR VPWR _03509_ sky130_fd_sc_hd__o2bb2ai_1
X_11529_ _02464_ _02465_ _02466_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__a21o_1
Xwire293 _03026_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__buf_4
X_18085_ _08880_ _08901_ _08931_ _08932_ VGND VGND VPWR VPWR _08934_ sky130_fd_sc_hd__o211a_1
X_15297_ _06110_ net944 net719 VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__and3_1
X_14317_ _05194_ _05196_ _05213_ _05215_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__o211ai_2
X_17036_ _07821_ net523 net554 VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__nand3_1
X_14248_ net771 net767 net656 net650 VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__nand4_2
XFILLER_98_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14179_ net210 net195 _05082_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__nand3_2
XFILLER_140_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_55_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18987_ net626 net718 _09873_ _09875_ VGND VGND VPWR VPWR _09878_ sky130_fd_sc_hd__a22oi_2
X_17938_ _08794_ _08769_ net795 _08795_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__o211a_1
XFILLER_78_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17869_ a_l\[12\] net473 VGND VGND VPWR VPWR _08729_ sky130_fd_sc_hd__nand2_1
XFILLER_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone172 net993 VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__clkbuf_16
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19608_ _09253_ _09308_ _00800_ _00801_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__o211ai_1
XFILLER_38_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19539_ _00631_ _00634_ net1002 _00680_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__a31o_1
XFILLER_62_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20314_ net793 net10 VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__and2_1
XFILLER_103_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap571 a_l\[11\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__clkbuf_8
Xmax_cap560 a_l\[13\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__buf_12
X_20245_ _01487_ _01488_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__and2b_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap582 net583 VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__buf_12
Xmax_cap593 net594 VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_8
XFILLER_67_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20176_ _01413_ _01414_ _09319_ _09362_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_103_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ net794 net1313 VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__and2_1
XFILLER_29_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11880_ _02816_ _02815_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_86_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ _01842_ _01846_ _01848_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10762_ p_hl\[21\] p_lh\[21\] VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__xor2_2
X_13550_ _04456_ _04436_ _04434_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12501_ net647 net644 net511 net508 VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__nand4_1
X_13481_ _04390_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__inv_2
XFILLER_139_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12432_ _03357_ _03360_ _03361_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a21bo_1
X_10693_ p_hl\[11\] p_lh\[11\] VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15220_ _06101_ _06105_ _06111_ _06112_ _06104_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__o221ai_2
XFILLER_138_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12363_ _03158_ _03286_ _03288_ _03276_ _03277_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__o2111ai_4
X_15151_ _06046_ _06047_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12294_ _09395_ _09679_ _03221_ _03222_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__o22ai_2
X_11314_ net691 net507 VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__nand2_2
XFILLER_107_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15082_ _05971_ _05976_ _05979_ _05975_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__o211ai_2
X_14102_ _04707_ _04923_ _04926_ _04922_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__a22o_2
XFILLER_141_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11245_ _02063_ _02068_ _02065_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__a21o_1
XFILLER_107_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14033_ _04934_ _04932_ _04937_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__a21o_1
X_18910_ net446 _09800_ _09798_ VGND VGND VPWR VPWR _09802_ sky130_fd_sc_hd__o21ai_1
XFILLER_122_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19890_ net568 net731 VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__nand2_1
X_11176_ _02116_ _02118_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__nand2_2
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18841_ _09313_ _09438_ _09587_ _09731_ _09590_ VGND VGND VPWR VPWR _09734_ sky130_fd_sc_hd__o2111ai_4
XFILLER_122_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15984_ net583 net541 VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__nand2_1
XFILLER_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18772_ _09660_ _09661_ VGND VGND VPWR VPWR _09662_ sky130_fd_sc_hd__nand2_1
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17723_ _08578_ _08579_ _08209_ _08375_ VGND VGND VPWR VPWR _08586_ sky130_fd_sc_hd__nand4_1
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14935_ _05823_ _05828_ net424 _05827_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_128_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17654_ _08511_ _08512_ _08514_ _08406_ VGND VGND VPWR VPWR _08518_ sky130_fd_sc_hd__o2bb2ai_4
X_14866_ _05756_ _05758_ _05759_ _05751_ _05749_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__o2111ai_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16605_ _07471_ _07472_ net629 net477 VGND VGND VPWR VPWR _07477_ sky130_fd_sc_hd__o211a_1
X_17585_ _08445_ _08352_ _08444_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__nand3_2
X_13817_ _04719_ _04721_ _04722_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__a21o_1
X_14797_ net806 _05695_ _05693_ _05692_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_141_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16536_ _07400_ _07405_ _07408_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__o21ai_1
X_13748_ _04647_ _04648_ _04625_ net287 VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__o211ai_4
X_19324_ _00497_ _00498_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__nand2_1
X_19255_ _10005_ _10154_ _10155_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__o21a_1
X_16467_ _07199_ _07204_ _07202_ VGND VGND VPWR VPWR _07340_ sky130_fd_sc_hd__a21boi_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18206_ _09188_ _09220_ _09049_ _09051_ VGND VGND VPWR VPWR _09053_ sky130_fd_sc_hd__o22a_1
X_13679_ _04503_ _04544_ _04542_ _04536_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_TAPCELL_ROW_42_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16398_ _07266_ _07267_ _07269_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__nand3_2
X_19186_ _10077_ _10078_ _09144_ _09362_ VGND VGND VPWR VPWR _10081_ sky130_fd_sc_hd__o2bb2a_1
X_15418_ net722 net640 net635 net726 VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__a22o_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18137_ net774 net971 VGND VGND VPWR VPWR _08985_ sky130_fd_sc_hd__nand2_1
X_15349_ _06151_ _06155_ _06179_ _06186_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__a2bb2oi_4
X_18068_ net790 net601 VGND VGND VPWR VPWR _08917_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17019_ net612 net608 _02588_ _07742_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__a31o_1
XFILLER_125_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20030_ _01197_ _01199_ _01254_ _01256_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__a22o_1
XFILLER_100_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20794_ clknet_leaf_6_clk _00434_ VGND VGND VPWR VPWR b_h\[0\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_81_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer223 net766 VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__buf_12
Xrebuffer201 a_h\[6\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer212 a_h\[4\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_20_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer256 a_l\[13\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer245 _09204_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__buf_1
Xrebuffer234 _09676_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__buf_6
Xrebuffer278 _01979_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__buf_1
XFILLER_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap390 _05337_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ _01952_ _01953_ net328 _01971_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20228_ _01369_ _01410_ _01416_ _01424_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__o211ai_2
XFILLER_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20159_ _01321_ _01332_ _01392_ _01393_ _01398_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__a41o_1
XFILLER_134_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12981_ _03904_ _03905_ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__nand2_1
X_11932_ _02707_ net511 net665 VGND VGND VPWR VPWR _02868_ sky130_fd_sc_hd__nand3_1
X_14720_ _05611_ _05619_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__and3_2
XFILLER_17_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11863_ net248 _02760_ _02796_ _02759_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__o211ai_1
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14651_ net761 net642 VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10814_ _01816_ _01822_ _01827_ _01821_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__and4bb_1
X_17370_ _08199_ _08200_ _08233_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__nand3_1
X_13602_ _04508_ _04510_ _09220_ _09428_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_45_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16321_ net620 net816 net496 net491 VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__and4_1
X_11794_ net1062 _02613_ _02608_ _02611_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__o22ai_4
X_14582_ _05480_ _05481_ _09308_ _09439_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__o2bb2ai_1
X_10745_ p_hl\[19\] p_lh\[19\] VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__xor2_1
X_13533_ _04440_ _04441_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__nand2_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16252_ _07091_ _06989_ _07124_ _07125_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__o211ai_4
X_10676_ p_hl\[8\] p_lh\[8\] VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__nand2_1
X_13464_ _04372_ _04374_ _04265_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a21o_1
X_19040_ _09816_ _09930_ VGND VGND VPWR VPWR _09931_ sky130_fd_sc_hd__nand2_4
X_16183_ _06939_ _06944_ _06946_ _07051_ _07052_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__o2111a_1
X_12415_ net692 net687 net483 net481 _03178_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__a41o_1
X_13395_ _04266_ _04267_ _04302_ _04303_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__nand4_1
X_15203_ net730 net651 VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__nand2_1
X_12346_ net633 net526 VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__nand2_1
XFILLER_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15134_ _06029_ _06022_ _06017_ _06027_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__o211ai_2
XFILLER_142_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12277_ _03061_ _03066_ _03201_ _03202_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__nand4_2
X_19942_ _01087_ _01163_ _01164_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__nand3_2
X_15065_ _05916_ _05918_ _05960_ _05961_ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__nand4_1
X_11228_ net664 net539 VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__nand2_2
X_19873_ _01037_ _01088_ _01089_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__nand3_1
X_14016_ net746 net689 VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11159_ _02099_ _02101_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__nand2_1
XFILLER_122_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18824_ _09714_ _09711_ _09710_ VGND VGND VPWR VPWR _09717_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_52_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_143_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15967_ _06842_ _06843_ _06844_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__a21boi_1
X_18755_ _09640_ _09641_ VGND VGND VPWR VPWR _09643_ sky130_fd_sc_hd__nand2_1
XFILLER_49_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15898_ net613 net515 _06774_ _06775_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__a22oi_2
X_17706_ net1054 net488 _08564_ _08567_ VGND VGND VPWR VPWR _08569_ sky130_fd_sc_hd__a22o_1
X_18686_ _09399_ _09400_ _09325_ _09421_ VGND VGND VPWR VPWR _09568_ sky130_fd_sc_hd__a31oi_2
X_14918_ _05812_ _05813_ net761 net636 VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__nand4_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17637_ _08398_ _08489_ _08498_ _08499_ VGND VGND VPWR VPWR _08501_ sky130_fd_sc_hd__o211a_1
XFILLER_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14849_ _05669_ _05746_ _05747_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__nand3_4
XFILLER_90_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17568_ _09253_ _09275_ _02589_ _08321_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__o31a_1
X_19307_ net298 _00452_ _00476_ _00478_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__o2bb2ai_2
X_16519_ net876 net522 VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__nand2_2
X_17499_ _08362_ _08363_ _08364_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19238_ _10117_ _10119_ _10132_ VGND VGND VPWR VPWR _10138_ sky130_fd_sc_hd__o21ai_2
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_19169_ _10059_ _10058_ _10032_ VGND VGND VPWR VPWR _10063_ sky130_fd_sc_hd__a21o_1
XFILLER_145_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20013_ _01104_ _01098_ _01238_ _01235_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__o22ai_2
XFILLER_100_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20777_ clknet_leaf_59_clk _00417_ VGND VGND VPWR VPWR a_h\[15\] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10530_ net795 net1202 VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__and2_1
X_10461_ term_mid\[45\] term_high\[45\] _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_98_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ _03130_ _03132_ _09471_ _09613_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_89_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10392_ term_mid\[36\] term_high\[36\] VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__xor2_1
X_13180_ _04100_ _04101_ _04078_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__a21o_1
X_12131_ _03045_ _03046_ _03062_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__o21ai_2
X_12062_ _02899_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nand2_2
Xhold490 mid_sum\[8\] VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
X_11013_ net691 net534 VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__and2_1
XFILLER_104_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16870_ net612 net608 net485 net479 VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__nand4_2
X_15821_ _06696_ _06697_ _06692_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__a21oi_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _06630_ net955 VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__nand2_2
X_12964_ net976 net1112 VGND VGND VPWR VPWR _03891_ sky130_fd_sc_hd__nand2_1
X_18540_ net630 net732 VGND VGND VPWR VPWR _09409_ sky130_fd_sc_hd__nand2_1
XFILLER_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11915_ _02848_ _02825_ _02847_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__nand3_1
X_18471_ net604 net759 net754 net887 VGND VGND VPWR VPWR _09333_ sky130_fd_sc_hd__a22oi_4
X_14703_ net723 net685 VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_107_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _06554_ _06556_ _06562_ _06557_ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__o211a_1
X_17422_ _08210_ _08286_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__nand2_1
XFILLER_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12895_ net976 net885 VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__nand2_1
X_11846_ _02780_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__nand2_1
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14634_ _05534_ _05533_ _05532_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__and3_1
X_11777_ _02703_ _02710_ _02711_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__nand3_2
X_17353_ _08043_ _08212_ _08213_ VGND VGND VPWR VPWR _08220_ sky130_fd_sc_hd__nand3_4
X_14565_ net727 net690 VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__nand2_4
X_16304_ net161 _07170_ _07174_ VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__a21o_1
X_17284_ _08148_ _08150_ VGND VGND VPWR VPWR _08152_ sky130_fd_sc_hd__nand2_1
X_10728_ _01756_ _01758_ net468 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a21oi_1
X_13516_ net433 _04420_ _04410_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__o21ai_2
X_16235_ net950 net515 VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__nand2_1
X_14496_ _05266_ _05397_ _05398_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__nand3_4
X_19023_ net457 _06985_ _09907_ _09910_ VGND VGND VPWR VPWR _09914_ sky130_fd_sc_hd__o211a_1
Xclkload35 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinv_4
Xclkload24 clknet_leaf_41_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_6
Xclkload13 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_4
X_10659_ _01698_ _01699_ _01700_ net797 VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__a31o_1
X_13447_ _04355_ _04356_ _04346_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__nand3_2
X_16166_ _07022_ _07023_ _07037_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__nand3_1
XFILLER_127_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload46 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__inv_8
X_13378_ _04286_ _04288_ _09155_ _09428_ VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_11_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16097_ _06968_ _06969_ _06971_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__nand3_1
X_12329_ net653 net647 net511 net508 VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__and4_1
X_15117_ net719 a_h\[8\] _06008_ _06011_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__a22oi_2
XFILLER_142_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19925_ _01142_ _01143_ _01145_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__nand3_1
X_15048_ net719 a_h\[7\] _05943_ _05944_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__a22o_1
XFILLER_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19856_ net603 net717 _00864_ _00862_ VGND VGND VPWR VPWR _01073_ sky130_fd_sc_hd__a31o_1
X_16999_ _07863_ _07865_ _07864_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__nand3_2
XFILLER_96_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18807_ _09688_ _09692_ _09694_ VGND VGND VPWR VPWR _09700_ sky130_fd_sc_hd__and3_1
X_19787_ _00888_ _00889_ net407 _00995_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__a31oi_2
X_18738_ _09595_ _09621_ _09623_ VGND VGND VPWR VPWR _09625_ sky130_fd_sc_hd__and3_1
X_20700_ clknet_leaf_39_clk _00340_ VGND VGND VPWR VPWR p_lh\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18669_ _09544_ _09546_ net630 net729 VGND VGND VPWR VPWR _09550_ sky130_fd_sc_hd__nand4_1
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20631_ clknet_leaf_50_clk _00271_ VGND VGND VPWR VPWR p_ll_pipe\[29\] sky130_fd_sc_hd__dfxtp_1
X_20562_ clknet_leaf_17_clk _00202_ VGND VGND VPWR VPWR mid_sum\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload7 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload7/X sky130_fd_sc_hd__clkbuf_4
X_20493_ clknet_leaf_27_clk _00133_ VGND VGND VPWR VPWR term_mid\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_286 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11700_ net462 _02633_ _02632_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__o21ai_1
X_12680_ _03502_ _03589_ _03591_ _03594_ _03500_ VGND VGND VPWR VPWR _03610_ sky130_fd_sc_hd__a32oi_1
XFILLER_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11631_ _02565_ _02567_ _02441_ net796 VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_120_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11562_ _02498_ _02499_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__nand2_2
XFILLER_24_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14350_ _05249_ _05252_ _04837_ _05087_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__o2bb2ai_2
X_10513_ term_high\[56\] term_high\[57\] term_high\[58\] VGND VGND VPWR VPWR _01664_
+ sky130_fd_sc_hd__and3_1
X_13301_ _04184_ _04188_ a_h\[0\] net757 VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o211ai_4
X_11493_ _02430_ _02432_ _02244_ _02245_ VGND VGND VPWR VPWR _02433_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14281_ _05144_ _05177_ _05178_ _05032_ _05006_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a32oi_1
X_10444_ term_mid\[42\] term_high\[42\] _01608_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__a21bo_1
X_16020_ net624 net502 VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__nand2_1
X_13232_ net784 net704 net700 net787 VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__a22o_1
X_10375_ _01417_ _01460_ net796 VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13163_ _04070_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__or2_1
X_12114_ _02837_ _02838_ _02834_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__a21oi_4
XFILLER_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17971_ _08819_ _08821_ net627 net779 VGND VGND VPWR VPWR _08823_ sky130_fd_sc_hd__nand4_1
X_13094_ _04017_ _04018_ _09493_ _09679_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__o2bb2ai_2
X_19710_ net1079 net574 b_l\[10\] VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__nand3_2
XFILLER_120_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16922_ _07780_ _07786_ VGND VGND VPWR VPWR _07792_ sky130_fd_sc_hd__nand2_1
X_12045_ _02864_ _02976_ _02978_ _02862_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__o2bb2ai_1
X_16853_ _07721_ _07723_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__nand2_1
XFILLER_93_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19641_ _00837_ _00839_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__nand2_1
X_15804_ net607 net602 net531 net527 VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__nand4_2
XFILLER_1_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19572_ net367 _00756_ _00760_ net406 VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__o211a_1
X_16784_ _07649_ _07650_ _07637_ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__nand3_2
X_18523_ _09380_ _09382_ _09364_ VGND VGND VPWR VPWR _09390_ sky130_fd_sc_hd__a21o_1
XFILLER_1_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13996_ _04896_ _04898_ _09155_ _09493_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__o2bb2ai_2
X_15735_ _06598_ _06611_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_105_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12947_ _03870_ _03874_ _03873_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__o21a_2
XFILLER_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15666_ _06530_ _06532_ _06542_ _06544_ net309 VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__o2111ai_1
X_18454_ _09312_ _09314_ net153 VGND VGND VPWR VPWR _09315_ sky130_fd_sc_hd__a21oi_4
X_12878_ _03507_ net633 VGND VGND VPWR VPWR _03806_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11829_ net712 net475 _02763_ _02765_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__a22oi_2
X_17405_ _08017_ _08019_ _08158_ VGND VGND VPWR VPWR _08272_ sky130_fd_sc_hd__o21ai_1
X_18385_ net791 net782 net584 net573 VGND VGND VPWR VPWR _09239_ sky130_fd_sc_hd__nand4_2
XFILLER_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14617_ _05506_ _05507_ _05514_ _05516_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_16_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15597_ _06476_ _06477_ VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__nand2_4
X_17336_ _08045_ _08046_ _08074_ _08077_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__o22ai_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14548_ _05271_ _05446_ net761 net649 _05445_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__o2111ai_4
X_17267_ _08125_ _08124_ _08082_ _08079_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__a22oi_1
X_14479_ _05024_ _05221_ _05222_ _05227_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__a31o_1
XFILLER_134_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16218_ _06980_ _06986_ _06982_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__a21oi_1
X_17198_ _08064_ _08061_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__nand2_1
X_19006_ net369 _09890_ VGND VGND VPWR VPWR _09897_ sky130_fd_sc_hd__nand2_1
X_16149_ _07022_ _07023_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19908_ net580 net574 net1043 net1099 VGND VGND VPWR VPWR _01129_ sky130_fd_sc_hd__nand4_1
XFILLER_110_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19839_ _01050_ _01052_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__nor2_2
XFILLER_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20614_ clknet_leaf_41_clk _00254_ VGND VGND VPWR VPWR p_ll_pipe\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20545_ clknet_leaf_43_clk net229 VGND VGND VPWR VPWR mid_sum\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20476_ clknet_leaf_43_clk _00116_ VGND VGND VPWR VPWR term_mid\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_122_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13850_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__inv_2
X_10993_ _01882_ _01902_ _01938_ _01901_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_122_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12801_ _03672_ b_h\[8\] net645 VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__nand3_1
X_13781_ _04687_ _04562_ _04681_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__nand3_2
X_15520_ net627 net540 net532 net631 VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__a22o_1
X_12732_ _03659_ _03523_ _03658_ VGND VGND VPWR VPWR _03662_ sky130_fd_sc_hd__nand3_2
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15451_ net155 _06333_ _06332_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__o21ai_1
X_12663_ _03593_ _03501_ _03592_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__nand3_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ net667 net662 net1125 VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__and3_1
X_11614_ _02545_ _02550_ _02447_ _02551_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_100_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _09016_ _09017_ VGND VGND VPWR VPWR _09018_ sky130_fd_sc_hd__nand2_1
X_12594_ _03514_ _03518_ _03517_ VGND VGND VPWR VPWR _03525_ sky130_fd_sc_hd__o21ai_1
X_15382_ _06233_ _06271_ _06272_ _06273_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__nand4_1
XFILLER_128_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11545_ net664 net526 net520 net672 VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__a22o_1
X_17121_ _07831_ _07837_ _07940_ _07943_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__nand4_2
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14333_ _05229_ _05231_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__nand2_1
Xmax_cap208 _07414_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_2
X_11476_ _02411_ _02413_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__nand2_1
X_17052_ net578 net503 VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__and2_1
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14264_ net454 _05166_ _05156_ _05167_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__o211ai_4
X_10427_ _01595_ net443 net796 VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_133_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16003_ net572 net521 VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__nand2_1
X_13215_ net1088 net784 VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__and2_2
Xmax_cap219 _08948_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__buf_6
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14195_ _05097_ _04960_ _05095_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__nand3_1
X_13146_ _04068_ _04031_ net793 _04069_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__o211a_1
X_10358_ _01161_ _01300_ _01289_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__o21ai_1
X_17954_ net796 _08808_ _08809_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__nor3_1
X_13077_ net641 net1112 VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__nand2_1
X_10289_ term_low\[20\] term_mid\[20\] _00471_ _00547_ VGND VGND VPWR VPWR _00569_
+ sky130_fd_sc_hd__o211ai_2
X_12028_ _02959_ _02963_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__and2_1
X_16905_ _07771_ _07772_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17885_ _08737_ _08740_ _08742_ _08739_ VGND VGND VPWR VPWR _08745_ sky130_fd_sc_hd__o211ai_1
XFILLER_66_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16836_ _07473_ _07474_ _07483_ _07487_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__a22o_1
X_19624_ _00817_ _00819_ _00820_ _00609_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__o2bb2ai_4
X_16767_ _07527_ _07534_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__nand2_1
X_19555_ _00746_ _00748_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__nand2_1
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13979_ _09220_ _09460_ _04876_ _04878_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__o22a_2
X_15718_ _06518_ _06522_ _06523_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__a21oi_1
X_18506_ net791 net569 VGND VGND VPWR VPWR _09371_ sky130_fd_sc_hd__nand2_2
X_19486_ _00643_ _00645_ _00670_ _00672_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16698_ _07560_ _07563_ _07565_ _07450_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__o211ai_1
X_18437_ _09227_ _09293_ _09294_ VGND VGND VPWR VPWR _09296_ sky130_fd_sc_hd__nand3_4
XFILLER_34_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15649_ _09188_ _09199_ _06440_ _06517_ _06524_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_32_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18368_ _09114_ _09122_ _09123_ _09127_ VGND VGND VPWR VPWR _09221_ sky130_fd_sc_hd__a31o_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18299_ _09063_ _09064_ _09061_ VGND VGND VPWR VPWR _09146_ sky130_fd_sc_hd__a21oi_1
X_17319_ _09231_ _09668_ _08180_ _08181_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__o22ai_2
X_20330_ net793 net23 VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__and2_1
XFILLER_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap720 b_l\[14\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__buf_6
Xmax_cap731 b_l\[11\] VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__buf_6
X_20261_ _01503_ _01504_ net557 b_l\[15\] VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__and4b_1
Xmax_cap753 net755 VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__buf_12
XFILLER_89_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap775 net776 VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__buf_12
Xmax_cap797 net65 VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__buf_12
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20192_ _01430_ _01431_ _01426_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__and3_1
Xmax_cap786 b_l\[1\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__buf_12
XFILLER_130_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11330_ _02266_ _02267_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__nand2_1
X_20528_ clknet_leaf_47_clk _00168_ VGND VGND VPWR VPWR term_low\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20459_ clknet_leaf_14_clk _00099_ VGND VGND VPWR VPWR term_high\[51\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11261_ _02199_ net361 _02201_ net464 VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o2bb2a_1
X_11192_ _02053_ _01984_ _02052_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_115_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13000_ _03925_ _03926_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__nand2_1
X_10212_ a_h\[11\] VGND VGND VPWR VPWR _09493_ sky130_fd_sc_hd__inv_6
XFILLER_121_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14951_ _05845_ _05846_ _05849_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__nand3_4
X_17670_ _08529_ _08530_ _08531_ VGND VGND VPWR VPWR _08534_ sky130_fd_sc_hd__nand3_2
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13902_ _04774_ _04776_ _04801_ _04803_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nand4_1
X_14882_ _05667_ _05769_ _05770_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__a21boi_2
X_16621_ _07390_ net453 VGND VGND VPWR VPWR _07493_ sky130_fd_sc_hd__nor2_1
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13833_ _04736_ _04737_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__nor2_2
X_16552_ _02588_ net848 _07219_ _07212_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__a22o_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19340_ _00499_ _00506_ _10091_ _10093_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__o211ai_2
X_10976_ net691 net686 net545 net538 VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__nand4_2
X_13764_ _04488_ _04498_ _04500_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15503_ _06364_ _06382_ _06383_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__o21a_1
XFILLER_15_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16483_ a_l\[7\] net590 net513 net506 VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__nand4_1
X_12715_ _09635_ _03639_ _03635_ _03642_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__o211ai_1
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13695_ _04596_ _04597_ _04591_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__a21o_1
XFILLER_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19271_ _09220_ _09319_ _10042_ _10170_ _10168_ VGND VGND VPWR VPWR _10173_ sky130_fd_sc_hd__o221ai_1
X_12646_ _03504_ _03570_ _03573_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__and3_1
X_18222_ _09066_ _09068_ _09155_ _09231_ VGND VGND VPWR VPWR _09069_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15434_ _06283_ _06287_ _06324_ _06325_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ _08963_ _08997_ _08998_ VGND VGND VPWR VPWR _09001_ sky130_fd_sc_hd__nand3_2
X_15365_ net156 _06255_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__nor2_1
X_17104_ net451 _07968_ _07966_ VGND VGND VPWR VPWR _07973_ sky130_fd_sc_hd__o21ai_4
X_12577_ net644 net1036 net964 net509 VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__nand4_1
X_14316_ _05199_ _05214_ _05213_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__o21a_1
Xwire283 _06815_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_2
Xwire261 _06816_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_2
X_11528_ _02464_ _02465_ _02466_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__a21oi_2
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18084_ _08930_ _08913_ _08902_ _08881_ VGND VGND VPWR VPWR _08933_ sky130_fd_sc_hd__a22oi_1
Xwire272 _00892_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_2
X_15296_ _06188_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__nor2_1
X_11459_ net692 net687 net1018 net507 VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__nand4_1
X_17035_ _07392_ net516 net1004 VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__nand3_1
X_14247_ _05148_ _05149_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__nand2_2
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14178_ _05037_ _05039_ _05077_ _05078_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_55_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _04011_ _04051_ _04008_ _04009_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__nand4b_1
XTAP_TAPCELL_ROW_55_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _09873_ _09875_ net1128 net718 VGND VGND VPWR VPWR _09877_ sky130_fd_sc_hd__and4_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17937_ _08793_ _08792_ VGND VGND VPWR VPWR _08795_ sky130_fd_sc_hd__nand2_1
XFILLER_93_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17868_ _08726_ _08727_ VGND VGND VPWR VPWR _08728_ sky130_fd_sc_hd__nand2_1
XFILLER_39_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16819_ _07680_ _07686_ _07685_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__o21ai_1
XFILLER_53_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19607_ _00800_ _00801_ _00802_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__a21o_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17799_ _08520_ _08590_ _08605_ VGND VGND VPWR VPWR _08661_ sky130_fd_sc_hd__o21ai_1
X_19538_ _00631_ _00634_ _00682_ _00680_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__a31oi_2
X_19469_ _09264_ _09286_ _00654_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__o21ai_2
XFILLER_61_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20313_ net793 net9 VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__and2_1
XFILLER_131_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap572 net578 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__buf_8
Xmax_cap561 net566 VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_12
Xmax_cap550 a_l\[15\] VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__buf_8
X_20244_ _01488_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__inv_2
XFILLER_143_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap594 a_l\[7\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_8
XFILLER_89_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20175_ _01411_ _01412_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__nand2_1
XFILLER_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10830_ _01842_ _01846_ net795 VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__o21ai_1
X_10761_ net442 _01782_ _01784_ _01788_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__o31a_1
X_12500_ net645 net508 VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__nand2_2
X_13480_ _04327_ net1125 net963 net714 _04328_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__a41o_1
X_10692_ _01725_ _01727_ _01729_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12431_ _03225_ _03228_ _03357_ _03360_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__nand4_1
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12362_ _03163_ _03291_ _03292_ _03293_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__nand4_4
X_15150_ _06004_ _06044_ _06045_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__nand3b_4
XFILLER_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12293_ _09395_ _09679_ _03221_ _03222_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__o22a_1
X_11313_ net706 net501 VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__nand2_1
X_15081_ _09384_ _09428_ _05784_ _05787_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__o31a_1
X_14101_ _05001_ _04971_ _04999_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_130_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11244_ _02153_ _02182_ _02183_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__nand3_4
XFILLER_106_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14032_ _04934_ _04932_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__a21oi_1
X_11175_ _02114_ _02115_ _02038_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__nand3_1
XFILLER_121_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18840_ _09437_ _09584_ _09728_ VGND VGND VPWR VPWR _09733_ sky130_fd_sc_hd__or3_1
XFILLER_121_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15983_ _06756_ _06759_ _06762_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__o21a_1
X_18771_ net792 net1064 net564 net560 VGND VGND VPWR VPWR _09661_ sky130_fd_sc_hd__nand4_4
X_17722_ _08579_ _08377_ VGND VGND VPWR VPWR _08585_ sky130_fd_sc_hd__nand2_1
X_14934_ _05717_ _05831_ _05830_ _05829_ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_145_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _08511_ _08512_ _08515_ VGND VGND VPWR VPWR _08517_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_50_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16604_ net629 net477 _07471_ _07472_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__a211oi_1
XPHY_EDGE_ROW_121_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14865_ _05752_ _05762_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__nand2_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17584_ _08445_ _08352_ _08444_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__and3_1
X_13816_ _04719_ _04721_ _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__a21oi_1
X_14796_ net745 _05573_ net662 net806 VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__a31o_1
XFILLER_16_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10959_ _01883_ _01884_ _01897_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__o21a_1
X_16535_ _07404_ _07403_ _07370_ VGND VGND VPWR VPWR _07408_ sky130_fd_sc_hd__nand3_4
X_13747_ _04587_ _04650_ _04651_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__nand3_4
X_19323_ net588 net744 net738 net592 VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__a22oi_4
X_16466_ _07199_ net420 _07202_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__a21bo_1
X_19254_ _10005_ _10154_ net797 VGND VGND VPWR VPWR _10155_ sky130_fd_sc_hd__a21oi_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18205_ net774 net610 net769 net605 VGND VGND VPWR VPWR _09052_ sky130_fd_sc_hd__nand4_2
X_13678_ _04505_ _04537_ _04538_ _04503_ _04544_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__a32oi_4
X_15417_ _06250_ _06289_ _06296_ VGND VGND VPWR VPWR _06309_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_42_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16397_ _07270_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__inv_2
XFILLER_129_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12629_ _03548_ _03557_ _03549_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__and3_1
X_19185_ _05044_ _06521_ net621 net718 _10078_ VGND VGND VPWR VPWR _10080_ sky130_fd_sc_hd__o2111ai_4
XPHY_EDGE_ROW_130_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18136_ net615 net769 VGND VGND VPWR VPWR _08984_ sky130_fd_sc_hd__nand2_1
X_15348_ _09362_ _09482_ _06149_ _06152_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__o31a_1
X_18067_ net779 net610 VGND VGND VPWR VPWR _08916_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15279_ _06168_ _06170_ _06159_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__a21oi_1
X_17018_ _09188_ _09679_ VGND VGND VPWR VPWR _07887_ sky130_fd_sc_hd__nor2_1
XFILLER_113_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18969_ _09722_ _09858_ _09726_ _09856_ VGND VGND VPWR VPWR _09861_ sky130_fd_sc_hd__and4_1
XFILLER_100_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20793_ clknet_leaf_8_clk _00433_ VGND VGND VPWR VPWR a_l\[15\] sky130_fd_sc_hd__dfxtp_4
XFILLER_35_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer213 net1009 VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_20_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer224 _02579_ VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer246 b_l\[12\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__buf_2
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer279 net711 VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_112_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20227_ _01411_ _01412_ _01416_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20158_ _01357_ _01395_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__nand2_1
XFILLER_134_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12980_ net634 net858 net824 net1049 VGND VGND VPWR VPWR _03907_ sky130_fd_sc_hd__a22oi_1
X_20089_ _01321_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__nand2_1
X_11931_ _02862_ net508 net672 VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__nand3_1
XFILLER_84_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11862_ _02761_ _02795_ VGND VGND VPWR VPWR _02799_ sky130_fd_sc_hd__nand2_1
XFILLER_72_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14650_ _05463_ _05550_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _01808_ _01818_ _01821_ _01827_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__and4b_1
X_13601_ _04402_ _04507_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nand2_1
X_14581_ _09308_ _09439_ _05480_ _05481_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__o211ai_1
X_16320_ _07191_ _07192_ VGND VGND VPWR VPWR _07194_ sky130_fd_sc_hd__nand2_1
X_11793_ _02728_ _02729_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__nand2_1
X_13532_ net757 net751 net705 net701 VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__nand4_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10744_ _01767_ _01771_ _01773_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__o21a_1
XFILLER_13_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16251_ _06989_ _07091_ _07125_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__o21ai_2
X_10675_ _09537_ _09548_ _01709_ _01711_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__o211ai_2
X_13463_ _04320_ _04368_ _04369_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__nand3_2
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16182_ _06841_ _06941_ _06949_ _07052_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__a22oi_2
XFILLER_127_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12414_ _03170_ _03213_ _03343_ _03344_ _03169_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__o2111ai_4
X_13394_ _04302_ _04303_ _04268_ VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__a21o_1
X_15202_ net730 net651 VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__and2_1
XFILLER_126_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12345_ net644 net518 VGND VGND VPWR VPWR _03278_ sky130_fd_sc_hd__nand2_1
X_15133_ _05930_ _05934_ _06022_ _06029_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_142_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12276_ _03202_ _03204_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__nand2_1
X_19941_ _01163_ _01164_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__nand2_1
X_15064_ _05918_ _05960_ _05961_ VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand3_1
X_11227_ _02166_ _02167_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__nand2_2
X_19872_ _01035_ _01003_ _01034_ _01039_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__a31o_1
X_14015_ _04734_ _04735_ _04732_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_147_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11158_ _02062_ _02094_ _02096_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__nand3_2
XFILLER_95_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18823_ _09715_ _09713_ _09712_ VGND VGND VPWR VPWR _09716_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_52_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_143_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11089_ _02029_ _02030_ _01999_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__a21oi_2
X_15966_ _06842_ _06843_ _09690_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__o21a_1
X_18754_ net1131 net581 net576 net775 VGND VGND VPWR VPWR _09642_ sky130_fd_sc_hd__a22oi_2
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15897_ net607 net583 net543 net521 VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__nand4_4
X_17705_ _09340_ _09646_ _08564_ _08567_ VGND VGND VPWR VPWR _08568_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18685_ _09529_ _09530_ _09562_ VGND VGND VPWR VPWR _09567_ sky130_fd_sc_hd__nand3_2
X_14917_ _05806_ _05808_ _05809_ _05674_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__a31o_1
X_17636_ _08498_ _08499_ VGND VGND VPWR VPWR _08500_ sky130_fd_sc_hd__nand2_1
X_14848_ _05744_ _05745_ _05670_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__a21oi_2
X_17567_ _09242_ _09679_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__nor2_1
X_16518_ net876 net544 net523 net572 VGND VGND VPWR VPWR _07391_ sky130_fd_sc_hd__a22oi_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14779_ _05552_ _05555_ _05553_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__a21oi_1
X_19306_ net298 _00452_ _00477_ _00479_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__nand4_2
X_17498_ _08264_ _08266_ _08265_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__a21boi_2
X_16449_ net812 net491 VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19237_ _10117_ _10119_ _10133_ VGND VGND VPWR VPWR _10136_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19168_ _10032_ _10058_ _10059_ VGND VGND VPWR VPWR _10062_ sky130_fd_sc_hd__nand3_2
XFILLER_145_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18119_ net781 net601 VGND VGND VPWR VPWR _08967_ sky130_fd_sc_hd__nand2_1
XFILLER_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19099_ _09983_ _09985_ _09976_ _09977_ VGND VGND VPWR VPWR _09990_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_6_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20012_ _01103_ _01099_ _01239_ _01237_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__a22oi_1
XFILLER_59_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ clknet_leaf_59_clk _00416_ VGND VGND VPWR VPWR a_h\[14\] sky130_fd_sc_hd__dfxtp_4
X_10460_ term_mid\[44\] term_high\[44\] term_mid\[45\] term_high\[45\] VGND VGND VPWR
+ VPWR _01623_ sky130_fd_sc_hd__a22o_1
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10391_ net470 _01563_ _01564_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__o21a_1
XFILLER_124_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12130_ _03047_ _03061_ _03062_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__nand3_2
XFILLER_145_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12061_ net637 net535 VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__nand2_4
Xhold480 mid_sum\[4\] VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold491 p_hh_pipe\[30\] VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11012_ _01918_ _01919_ _01922_ _01917_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a22oi_2
XFILLER_104_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15820_ _06696_ _06697_ net1127 net515 VGND VGND VPWR VPWR _06699_ sky130_fd_sc_hd__and4_1
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_125_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ net384 _06583_ _06626_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__o21ai_1
X_12963_ net659 net478 VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__and2_1
XFILLER_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11914_ _02846_ net399 VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__nand2_1
X_15682_ _06562_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__inv_2
XFILLER_73_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18470_ net604 net759 VGND VGND VPWR VPWR _09332_ sky130_fd_sc_hd__nand2_1
X_14702_ _05466_ _05602_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_107_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ net554 net550 net964 net969 VGND VGND VPWR VPWR _08287_ sky130_fd_sc_hd__nand4_4
XFILLER_61_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12894_ _09504_ _09646_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__nor2_1
X_14633_ _05532_ _05533_ _05534_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__a21oi_1
X_11845_ _02769_ _02778_ _02779_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__nand3b_2
X_11776_ _02706_ _02709_ _02704_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__a21o_1
X_17352_ _08042_ _08216_ _08215_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__nand3_2
X_14564_ net723 net690 VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__nand2_1
X_16303_ net161 _07170_ _07174_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__a21oi_2
X_17283_ _08145_ _08147_ _08150_ VGND VGND VPWR VPWR _08151_ sky130_fd_sc_hd__and3_1
X_10727_ _01756_ _01758_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__nand2_1
X_13515_ _09155_ _09449_ _04418_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__o21ai_1
X_14495_ _05377_ _05378_ _05387_ _05388_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__o2bb2ai_2
X_16234_ _07093_ _07106_ _07104_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__nand3_4
X_13446_ _04350_ _04354_ net434 VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__o21ai_4
XFILLER_9_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19022_ net592 net748 _09910_ _09911_ VGND VGND VPWR VPWR _09913_ sky130_fd_sc_hd__a22o_1
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10658_ _01699_ _01700_ _01698_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__a21oi_1
Xclkload14 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinv_1
Xclkload25 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_4
X_16165_ _07022_ _07023_ net1114 _07036_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__o2bb2ai_1
X_10589_ net793 net1302 VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__and2_1
Xclkload36 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__inv_12
Xclkload47 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinv_8
X_13377_ _04288_ net986 net777 VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_11_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16096_ _06968_ _06969_ _06970_ _06899_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__o2bb2ai_1
X_12328_ net647 net508 VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__nand2_4
X_15116_ _09362_ _06010_ _09460_ _06008_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__or4b_1
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ _03192_ _03182_ _03191_ VGND VGND VPWR VPWR _03193_ sky130_fd_sc_hd__and3_1
X_19924_ _01142_ _01143_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__a21o_1
X_15047_ net719 a_h\[7\] _05943_ _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__a22oi_2
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19855_ _01068_ _01071_ VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__nand2_1
X_16998_ _07861_ _07862_ _07866_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__nand3_2
X_18806_ _09692_ _09694_ VGND VGND VPWR VPWR _09699_ sky130_fd_sc_hd__nand2_1
X_19786_ _00888_ _00995_ _00889_ net407 VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__nand4_1
XFILLER_37_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15949_ net261 _06821_ _06823_ net262 VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__o211ai_1
XFILLER_110_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18737_ _09596_ _09597_ net335 _09619_ VGND VGND VPWR VPWR _09623_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18668_ _09544_ net729 net630 VGND VGND VPWR VPWR _09549_ sky130_fd_sc_hd__nand3_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17619_ net1093 a_l\[11\] net485 net479 VGND VGND VPWR VPWR _08483_ sky130_fd_sc_hd__nand4_1
X_18599_ _09470_ _09472_ VGND VGND VPWR VPWR _09473_ sky130_fd_sc_hd__nand2_2
XFILLER_51_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20630_ clknet_leaf_50_clk _00270_ VGND VGND VPWR VPWR p_ll_pipe\[28\] sky130_fd_sc_hd__dfxtp_1
X_20561_ clknet_leaf_17_clk _00201_ VGND VGND VPWR VPWR mid_sum\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkload8 clknet_leaf_57_clk VGND VGND VPWR VPWR clkload8/X sky130_fd_sc_hd__clkbuf_4
X_20492_ clknet_leaf_27_clk _00132_ VGND VGND VPWR VPWR term_mid\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11630_ _02565_ _02567_ _02441_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ net646 net546 net539 net652 VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__a22oi_4
XFILLER_70_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10512_ term_high\[56\] net1376 _01660_ net1358 VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__a31o_1
XFILLER_128_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13300_ a_h\[0\] net757 _04184_ _04188_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__a211o_1
XFILLER_7_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20759_ clknet_leaf_52_clk _00399_ VGND VGND VPWR VPWR p_ll\[29\] sky130_fd_sc_hd__dfxtp_1
X_11492_ _02337_ _02425_ _02426_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__nand3_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14280_ _05140_ _05142_ _05177_ _05178_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__nand4_4
X_10443_ term_mid\[43\] term_high\[43\] VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__xor2_1
X_13231_ net787 net784 net704 net700 VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__nand4_1
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10374_ _01417_ _01460_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__and2_1
XFILLER_108_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13162_ net225 _04084_ _04083_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__o21ai_2
X_12113_ _02837_ _02838_ _02834_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__a21o_1
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17970_ net627 net779 _08819_ _08821_ VGND VGND VPWR VPWR _08822_ sky130_fd_sc_hd__a22o_1
X_13093_ _03975_ _04015_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__nand2_2
X_12044_ net665 net658 net511 net508 VGND VGND VPWR VPWR _02979_ sky130_fd_sc_hd__nand4_1
X_16921_ _09275_ _09613_ _07671_ _07781_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__o22a_1
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16852_ _07722_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__inv_2
XFILLER_49_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19640_ _00726_ _00728_ _00835_ _00836_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__nand4_1
X_15803_ net607 net966 net531 net527 VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__and4_1
X_16783_ _07527_ _07534_ _07650_ VGND VGND VPWR VPWR _07654_ sky130_fd_sc_hd__nand3_1
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19571_ _00761_ _00763_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__nand2_1
X_15734_ _06613_ _06597_ _06612_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__nand3_4
X_18522_ _09237_ _09381_ _09380_ _09364_ VGND VGND VPWR VPWR _09389_ sky130_fd_sc_hd__o211ai_1
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_57_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_8
X_13995_ _04896_ _04898_ _04891_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__a21oi_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12946_ _03782_ _03784_ _03868_ _03867_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__o2bb2ai_1
X_15665_ _06542_ _06544_ VGND VGND VPWR VPWR _06546_ sky130_fd_sc_hd__nand2_2
X_18453_ _09305_ _09309_ _09205_ _09307_ VGND VGND VPWR VPWR _09314_ sky130_fd_sc_hd__o211ai_1
X_12877_ _03799_ _03800_ net674 net474 VGND VGND VPWR VPWR _03805_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_47_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11828_ net708 net706 net483 net481 VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__nand4_1
X_15596_ net616 net531 net527 net625 VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__a22oi_1
X_17404_ _08269_ _08270_ VGND VGND VPWR VPWR _08271_ sky130_fd_sc_hd__nand2_1
X_18384_ _09235_ _09236_ VGND VGND VPWR VPWR _09238_ sky130_fd_sc_hd__nand2_2
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14616_ _05513_ _05515_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_16_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _08115_ _08119_ _08193_ _08195_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__o211ai_1
X_14547_ _05447_ _05440_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__nand2_1
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11759_ _02602_ _02600_ _02590_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_60_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17266_ _08084_ _08086_ _08127_ _08129_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__o2bb2ai_2
X_14478_ _05217_ _05218_ _05023_ _05226_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__a31o_1
X_16217_ _09286_ _09581_ _06866_ _06981_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__o22a_1
X_17197_ _08053_ _08062_ _07903_ VGND VGND VPWR VPWR _08065_ sky130_fd_sc_hd__o21ai_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13429_ net772 net986 VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__nand2_1
X_19005_ _09877_ _09878_ _09895_ VGND VGND VPWR VPWR _09896_ sky130_fd_sc_hd__o21ai_2
X_16148_ _07023_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__inv_2
XFILLER_142_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16079_ _06876_ _06881_ _06879_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19907_ net580 net574 _05043_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__and3_1
XFILLER_96_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19838_ _01052_ _01050_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__nand2_4
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_28_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19769_ net797 _00977_ _00979_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_48_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20613_ clknet_leaf_41_clk _00253_ VGND VGND VPWR VPWR p_ll_pipe\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_61_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20544_ clknet_leaf_43_clk _00184_ VGND VGND VPWR VPWR mid_sum\[7\] sky130_fd_sc_hd__dfxtp_1
X_20475_ clknet_leaf_43_clk _00115_ VGND VGND VPWR VPWR term_mid\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_8
X_12800_ net634 net993 b_h\[8\] net1049 VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__a22oi_2
X_10992_ _01934_ _01936_ _01935_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__a21oi_2
X_13780_ _04681_ _04687_ _04558_ _04560_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_55_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12731_ _03659_ _03523_ _03658_ VGND VGND VPWR VPWR _03661_ sky130_fd_sc_hd__and3_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12662_ _03579_ _03587_ VGND VGND VPWR VPWR _03593_ sky130_fd_sc_hd__nand2_1
X_15450_ _06217_ _06340_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__nand2_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11613_ _02548_ _02549_ _02448_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__a21oi_2
XFILLER_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ net756 net750 net667 VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__nand3_1
X_17120_ _07830_ _07833_ _07946_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__a21oi_2
X_12593_ net353 _03516_ _03518_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15381_ _06227_ _06231_ _06273_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__o21a_1
XFILLER_129_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11544_ net664 net525 net1059 net671 VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__a22oi_4
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire432 _04666_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_2
X_14332_ _05233_ _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__nand2_1
Xwire410 _09928_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_1
X_11475_ _02407_ _02410_ _02408_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__and3_1
X_17051_ net1069 _07783_ net503 _07785_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__a31o_1
X_14263_ _05161_ _05163_ _05158_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__a21o_1
X_10426_ _01570_ _01591_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__a21o_2
X_16002_ _06877_ _06878_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__nand2_4
X_13214_ _09690_ net713 net791 VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__and3_1
Xwire498 net500 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_6
XFILLER_98_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14194_ _04955_ _04958_ _04957_ _05097_ _05095_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__a32o_1
X_13145_ _04031_ _04039_ _04067_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__o21bai_1
X_10357_ _01084_ _01095_ _01192_ _01203_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__or4_1
X_17953_ _08807_ _08799_ VGND VGND VPWR VPWR _08810_ sky130_fd_sc_hd__nand2_1
X_13076_ _09504_ _09668_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__nor2_1
X_10288_ term_low\[19\] term_mid\[19\] _00547_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12027_ _02960_ _02953_ _02809_ _02961_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o211ai_1
X_16904_ _07766_ _07770_ _07772_ VGND VGND VPWR VPWR _07774_ sky130_fd_sc_hd__nand3_2
XFILLER_25_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17884_ _08737_ _08740_ _08742_ _08739_ VGND VGND VPWR VPWR _08744_ sky130_fd_sc_hd__o211a_1
XFILLER_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19623_ _00607_ _00623_ _00609_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__a21oi_1
X_16835_ net629 net472 VGND VGND VPWR VPWR _07706_ sky130_fd_sc_hd__nand2_1
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16766_ _07524_ _07526_ _07528_ VGND VGND VPWR VPWR _07637_ sky130_fd_sc_hd__o21ai_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19554_ _00653_ _00744_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__nand2_4
X_13978_ _04879_ net670 net762 _04877_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__and4_4
X_16697_ _07564_ _07565_ _07450_ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__and3_1
X_15717_ _06518_ _06522_ _06523_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__a21o_1
XFILLER_80_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12929_ _03772_ _03855_ _03856_ VGND VGND VPWR VPWR _03857_ sky130_fd_sc_hd__nand3b_4
X_18505_ net782 net577 VGND VGND VPWR VPWR _09370_ sky130_fd_sc_hd__nand2_1
X_19485_ _00459_ _00663_ net833 _00661_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__o211ai_2
X_18436_ _09171_ _09226_ _09292_ VGND VGND VPWR VPWR _09295_ sky130_fd_sc_hd__nand3_4
X_15648_ net1120 net611 net531 net527 _06518_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_32_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15579_ _06433_ _06434_ _06447_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__o21a_1
X_18367_ net1082 net737 net847 _09218_ VGND VGND VPWR VPWR _09219_ sky130_fd_sc_hd__a31o_1
X_17318_ _09231_ _09668_ _08180_ _08181_ VGND VGND VPWR VPWR _08185_ sky130_fd_sc_hd__o22a_1
X_18298_ _09137_ _09143_ _09142_ VGND VGND VPWR VPWR _09145_ sky130_fd_sc_hd__o21ai_1
X_17249_ net342 _08116_ VGND VGND VPWR VPWR _08117_ sky130_fd_sc_hd__nand2_1
Xmax_cap710 net711 VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__buf_12
Xmax_cap721 b_l\[14\] VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__buf_8
X_20260_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__inv_2
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap732 b_l\[11\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__buf_6
Xmax_cap754 net755 VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkbuf_8
Xmax_cap743 net744 VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__buf_12
XFILLER_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap787 net789 VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__buf_8
X_20191_ _01431_ _01426_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__nand2_1
Xmax_cap765 b_l\[5\] VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__buf_12
Xmax_cap776 b_l\[3\] VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__buf_12
XFILLER_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_16_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_25_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20527_ clknet_leaf_47_clk _00167_ VGND VGND VPWR VPWR term_low\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20458_ clknet_leaf_14_clk _00098_ VGND VGND VPWR VPWR term_high\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11260_ _02108_ _02109_ net464 VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__a21oi_1
XFILLER_21_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11191_ _01984_ _02053_ _02051_ _02049_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_115_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10211_ net659 VGND VGND VPWR VPWR _09482_ sky130_fd_sc_hd__inv_8
X_20389_ clknet_leaf_41_clk _00029_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14950_ _05678_ _05690_ _05848_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__o21ai_2
XFILLER_87_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_34_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13901_ _04774_ _04801_ _04803_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__nand3_1
X_14881_ _05779_ _05780_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__nor2_1
X_16620_ _07260_ _07355_ _07360_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__o21ai_2
X_13832_ _04732_ _04734_ _04735_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__a21oi_1
X_16551_ _07220_ _07214_ _02589_ _06402_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__a211oi_2
XFILLER_62_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13763_ _04488_ _04498_ _04500_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__a21o_1
X_10975_ net686 net538 VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__nand2_4
X_12714_ _03640_ _03642_ _09482_ _09646_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__o2bb2ai_1
X_15502_ _06390_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__inv_2
X_16482_ net590 net506 VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__nand2_1
X_13694_ _02362_ _04134_ net777 net666 _04596_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_44_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19270_ _10166_ _10167_ _10170_ _10042_ VGND VGND VPWR VPWR _10172_ sky130_fd_sc_hd__o2bb2ai_1
X_12645_ _03574_ _03575_ _03503_ VGND VGND VPWR VPWR _03576_ sky130_fd_sc_hd__nand3_2
X_18221_ _09063_ _09064_ VGND VGND VPWR VPWR _09068_ sky130_fd_sc_hd__nand2_2
XPHY_EDGE_ROW_43_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15433_ _06322_ _06323_ _06316_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__a21o_1
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18152_ _08964_ _08995_ _08996_ VGND VGND VPWR VPWR _09000_ sky130_fd_sc_hd__nand3_2
X_12576_ net638 net509 VGND VGND VPWR VPWR _03507_ sky130_fd_sc_hd__nand2_1
X_15364_ _06255_ _06256_ net156 VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__o21ai_2
XFILLER_7_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11527_ _02392_ _02406_ _02412_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__o21ai_2
X_17103_ _09199_ _09668_ _07967_ _07968_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__o22a_1
X_18083_ _08930_ _08913_ VGND VGND VPWR VPWR _08932_ sky130_fd_sc_hd__nand2_2
X_14315_ _05199_ _05214_ _05213_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__o21ai_2
XFILLER_8_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17034_ net558 net554 net1023 net516 VGND VGND VPWR VPWR _07903_ sky130_fd_sc_hd__nand4_2
Xwire273 _00765_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__buf_1
X_15295_ _06127_ _06187_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__nor2_4
X_11458_ net692 net687 net1018 net507 VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__and4_1
X_14246_ net767 net656 net650 net771 VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__a22oi_1
X_10409_ _01578_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__nor2_1
X_11389_ _02321_ _02327_ _02329_ _02326_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__o211ai_1
XFILLER_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14177_ _05037_ _05039_ _05081_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__nand3_1
XFILLER_124_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _04011_ _04051_ _04008_ _04009_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__and4b_1
X_18985_ _09875_ net718 net1128 VGND VGND VPWR VPWR _09876_ sky130_fd_sc_hd__and3_1
X_17936_ _08788_ _08790_ _08770_ _08777_ VGND VGND VPWR VPWR _08794_ sky130_fd_sc_hd__o22ai_1
X_13059_ _03923_ _03978_ _03980_ _03977_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__a31o_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_94_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17867_ _08672_ _08684_ _08685_ _08725_ VGND VGND VPWR VPWR _08727_ sky130_fd_sc_hd__nand4b_2
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16818_ _07496_ _07682_ _07681_ _07678_ VGND VGND VPWR VPWR _07689_ sky130_fd_sc_hd__o211a_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19606_ _00800_ _00801_ _09253_ _09308_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__o2bb2ai_1
X_17798_ _08657_ _08659_ VGND VGND VPWR VPWR _08660_ sky130_fd_sc_hd__nand2_1
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19537_ _00726_ _00728_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__nand2_1
X_16749_ _07617_ _07592_ _07616_ VGND VGND VPWR VPWR _07620_ sky130_fd_sc_hd__nand3_2
XFILLER_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19468_ net896 net575 VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__and2_1
XFILLER_34_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18419_ _09144_ _09264_ net457 _06521_ _09274_ VGND VGND VPWR VPWR _09277_ sky130_fd_sc_hd__o221ai_4
XFILLER_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19399_ _00525_ _00527_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__nand2_1
XFILLER_147_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20312_ net793 net8 VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__and2_1
Xmax_cap540 net541 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_12
X_20243_ _01457_ _01486_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__or2_1
Xmax_cap551 net553 VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__buf_8
Xmax_cap562 net563 VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_12
Xmax_cap595 a_l\[7\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__buf_6
XFILLER_107_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap573 net578 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__buf_6
X_20174_ net727 net557 net724 net551 VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__nand4_1
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10760_ _01777_ _01778_ _01786_ net795 VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__o31a_1
XFILLER_52_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10691_ _01725_ _01727_ net794 VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12430_ _03360_ _03361_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__nand2_1
XFILLER_9_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12361_ _03144_ _03145_ _03163_ _03161_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__a31oi_2
X_14100_ _04971_ _04999_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__nand2_1
X_12292_ _09395_ _09679_ VGND VGND VPWR VPWR _03226_ sky130_fd_sc_hd__nor2_1
X_11312_ _02155_ _02160_ _02157_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__a21oi_1
X_15080_ _05785_ net690 net715 _05786_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_130_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11243_ _02181_ _02152_ _02180_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__nand3_2
X_14031_ _04932_ _04933_ _04918_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__a21oi_2
XFILLER_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11174_ _02114_ _02038_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__nand2_1
XFILLER_122_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15982_ _06756_ _06759_ _06762_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18770_ _09481_ _09658_ VGND VGND VPWR VPWR _09660_ sky130_fd_sc_hd__nand2_1
X_17721_ _08582_ _08581_ VGND VGND VPWR VPWR _08584_ sky130_fd_sc_hd__nand2_1
X_14933_ _05715_ _05719_ _05717_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_145_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17652_ _08392_ _08403_ _08404_ _08514_ VGND VGND VPWR VPWR _08516_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_50_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16603_ net629 net477 _07471_ _07472_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14864_ _05749_ _05751_ _05760_ _05761_ VGND VGND VPWR VPWR _05764_ sky130_fd_sc_hd__nand4_2
X_17583_ _08353_ _08446_ _08447_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__nand3_2
X_13815_ _09264_ _09406_ _04633_ _04635_ _04490_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__o32a_1
X_14795_ _05573_ net662 net745 VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__and3_1
X_10958_ _01882_ _01902_ _01904_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__a21oi_1
X_16534_ _07401_ _07402_ _07369_ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__nand3_1
XFILLER_50_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13746_ _04587_ _04651_ _04650_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__and3_1
XFILLER_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19322_ net588 net744 VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__nand2_1
X_16465_ _07271_ _07311_ _07336_ _07337_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__o211ai_2
XFILLER_92_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13677_ net1130 _04550_ _04584_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__o21ai_2
X_19253_ _10152_ _10153_ VGND VGND VPWR VPWR _10154_ sky130_fd_sc_hd__nand2_1
X_12628_ _03548_ _03549_ _03557_ VGND VGND VPWR VPWR _03559_ sky130_fd_sc_hd__a21o_1
X_18204_ net774 net610 net769 net605 VGND VGND VPWR VPWR _09051_ sky130_fd_sc_hd__and4_1
X_10889_ net794 net1219 VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__and2_1
X_15416_ net65 _06307_ _06308_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_42_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16396_ _07266_ _07267_ _07111_ _07268_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__o2bb2ai_4
X_19184_ _10078_ net718 net621 _10077_ VGND VGND VPWR VPWR _10079_ sky130_fd_sc_hd__and4_1
X_12559_ _03488_ _03489_ _03490_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a21oi_2
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18135_ net623 net764 VGND VGND VPWR VPWR _08983_ sky130_fd_sc_hd__nand2_1
X_15347_ _09384_ _09482_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__nor2_1
X_18066_ _08872_ _08869_ _08874_ VGND VGND VPWR VPWR _08915_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_57_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15278_ _06159_ _06168_ _06170_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__nand3_1
XFILLER_8_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17017_ _07869_ _07871_ VGND VGND VPWR VPWR _07886_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14229_ _05012_ _05126_ net746 net676 _05125_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__o2111ai_1
XFILLER_140_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18968_ _09726_ _09722_ _09858_ _09856_ VGND VGND VPWR VPWR _09860_ sky130_fd_sc_hd__a22oi_2
X_17919_ _08770_ net831 net795 VGND VGND VPWR VPWR _08778_ sky130_fd_sc_hd__o21ai_1
X_18899_ _09786_ _09787_ _09788_ VGND VGND VPWR VPWR _09791_ sky130_fd_sc_hd__a21o_1
XFILLER_82_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20792_ clknet_leaf_8_clk _00432_ VGND VGND VPWR VPWR a_l\[14\] sky130_fd_sc_hd__dfxtp_4
Xrebuffer214 net1009 VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_20_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer203 _05288_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_147_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer225 net500 VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_20_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer247 net1043 VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__buf_1
XFILLER_147_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer258 _05792_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer269 b_l\[1\] VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap381 _06885_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_112_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20226_ _09319_ _09384_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__nor2_1
Xmax_cap392 _04979_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_6
XFILLER_104_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20157_ _01321_ _01332_ _01392_ _01393_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__nand4_2
XFILLER_94_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11930_ _02863_ _02865_ net679 net501 VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__nand4_4
XFILLER_94_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20088_ _01252_ _01319_ _01320_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_127_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11861_ net248 _02760_ _02759_ _02795_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__o211ai_2
XFILLER_45_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _02724_ _02726_ net665 net518 VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand4_2
X_10812_ _01830_ _01831_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__nor2_1
XFILLER_72_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13600_ net768 net683 net675 net924 VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__a22oi_4
X_14580_ _05480_ _05481_ _05478_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_140_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _01771_ _01767_ net796 VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__a21oi_1
X_13531_ net757 net701 VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__nand2_1
X_16250_ _07108_ _07109_ _07120_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__a21o_1
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10674_ _01713_ _01714_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__nor2_1
X_13462_ _04320_ _04368_ _04369_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and3_1
X_15201_ _06091_ _06092_ _06095_ _06019_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__o2bb2ai_1
X_16181_ _07054_ _07055_ _07056_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__o21a_2
X_12413_ _03345_ _03342_ _03341_ VGND VGND VPWR VPWR _03346_ sky130_fd_sc_hd__nand3_4
X_13393_ _04302_ _04303_ _04268_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__a21bo_1
XFILLER_126_335 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12344_ _03254_ _03268_ _03269_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__nand3_1
X_15132_ _06019_ _06020_ _06018_ VGND VGND VPWR VPWR _06029_ sky130_fd_sc_hd__o21ai_2
X_19940_ _01157_ _01158_ _01097_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__a21o_1
X_15063_ _05955_ _05957_ _05920_ VGND VGND VPWR VPWR _05961_ sky130_fd_sc_hd__a21o_1
XFILLER_141_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12275_ _03061_ _03066_ _03201_ _03202_ VGND VGND VPWR VPWR _03209_ sky130_fd_sc_hd__a22o_1
X_14014_ _04732_ _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__nand2_1
X_11226_ net664 net965 net539 net671 VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__a22oi_1
X_19871_ net729 net725 _06984_ _01009_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__a31o_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ _02062_ _02094_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__nand2_1
X_18822_ _09562_ _09530_ _09527_ _09522_ VGND VGND VPWR VPWR _09715_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_52_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18753_ net768 net580 VGND VGND VPWR VPWR _09641_ sky130_fd_sc_hd__nand2_1
X_11088_ _02015_ _02017_ net403 _02025_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__o2bb2ai_1
X_15965_ _06570_ _06645_ _06730_ _06739_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__o31a_1
X_17704_ _08494_ _08565_ VGND VGND VPWR VPWR _08567_ sky130_fd_sc_hd__nand2_1
X_15896_ _06467_ _06772_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__nand2_2
X_18684_ _09529_ _09530_ _09562_ VGND VGND VPWR VPWR _09566_ sky130_fd_sc_hd__a21o_1
X_14916_ _05810_ _05805_ _05674_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__o21ai_2
X_17635_ _08496_ _08497_ VGND VGND VPWR VPWR _08499_ sky130_fd_sc_hd__nand2_1
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14847_ _05742_ _05740_ _05706_ _05707_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__o211ai_2
XFILLER_17_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17566_ _08299_ _08374_ _08425_ _08427_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_16_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16517_ net583 net516 VGND VGND VPWR VPWR _07390_ sky130_fd_sc_hd__nand2_2
X_14778_ _05552_ _05555_ _05553_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__a21o_1
X_19305_ _00463_ _00468_ _00470_ net1065 VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__o211ai_2
XFILLER_32_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17497_ _08248_ _08253_ _08359_ _08360_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__nand4_2
XFILLER_31_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13729_ net757 net752 net694 net689 _04631_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__a41o_1
X_16448_ _07191_ _07192_ _07190_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19236_ _10118_ _10120_ _10129_ _10131_ VGND VGND VPWR VPWR _10135_ sky130_fd_sc_hd__nand4_2
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16379_ _07240_ _07241_ _07251_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__a21o_1
X_19167_ _10058_ _10059_ VGND VGND VPWR VPWR _10060_ sky130_fd_sc_hd__nand2_1
X_18118_ net790 net594 VGND VGND VPWR VPWR _08966_ sky130_fd_sc_hd__nand2_1
XFILLER_145_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19098_ _09983_ _09985_ _09977_ VGND VGND VPWR VPWR _09989_ sky130_fd_sc_hd__o21ai_1
XFILLER_99_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18049_ _08895_ _08896_ VGND VGND VPWR VPWR _08898_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20011_ _01237_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__nand2_1
XFILLER_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_82_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20775_ clknet_leaf_0_clk _00415_ VGND VGND VPWR VPWR a_h\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10390_ _01563_ net470 net796 VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold481 p_hh\[15\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 p_hh_pipe\[29\] VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_12060_ _02987_ _02993_ _02992_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__o21ai_1
XFILLER_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11011_ _01918_ _01919_ _01922_ _01917_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_8_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20209_ _01343_ _01344_ _01402_ _01403_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__and4b_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold492 mid_sum\[5\] VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _06586_ _06618_ _06619_ _06584_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__a31oi_4
X_12962_ _09471_ _09679_ _03881_ _03882_ VGND VGND VPWR VPWR _03889_ sky130_fd_sc_hd__o211ai_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11913_ net399 _02843_ _02845_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__nand3b_1
X_15681_ _06496_ _06561_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__nand2_1
X_12893_ _03744_ _03749_ _03747_ VGND VGND VPWR VPWR _03821_ sky130_fd_sc_hd__a21oi_1
X_14701_ net727 net685 VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__nand2_1
X_11844_ _02776_ _02777_ _02769_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_107_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17420_ net550 net964 VGND VGND VPWR VPWR _08286_ sky130_fd_sc_hd__nand2_1
X_14632_ _05406_ _05263_ _05408_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_107_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11775_ _09439_ _09613_ _02650_ _02707_ _02706_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__o221ai_1
X_17351_ _08216_ _08042_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__nand2_1
XFILLER_60_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14563_ _05463_ _05464_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__nand2_1
X_16302_ _07045_ _07173_ _07170_ net161 VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__o211ai_4
X_17282_ _08149_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__inv_2
X_10726_ p_hl\[15\] p_lh\[15\] _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__a21oi_4
X_13514_ _04415_ _04417_ _04419_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__a21oi_2
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14494_ _05389_ _05390_ _05377_ _05378_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__o211ai_2
X_16233_ _06982_ _07092_ _07103_ _07105_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__o22ai_4
X_10657_ p_hl\[5\] p_lh\[5\] VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__or2_1
X_13445_ _09155_ _09439_ _02082_ _04134_ _04351_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__o221ai_2
X_19021_ _09910_ _09911_ _09907_ VGND VGND VPWR VPWR _09912_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload26 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_16
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload15 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__clkinv_8
Xclkload37 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__inv_16
X_16164_ net1114 _07036_ _07022_ _07023_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__o211ai_2
X_10588_ net793 net1257 VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__and2_1
Xclkload48 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_8
X_13376_ net787 net784 net932 net675 VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_11_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16095_ _06897_ _06902_ _06899_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__a21oi_2
X_12327_ _03131_ _03258_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__nand2_2
X_15115_ _06008_ _06011_ net719 a_h\[8\] VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__and4_1
XFILLER_114_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12258_ net682 net489 _03186_ _03187_ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__a22o_1
X_19923_ _01009_ _01011_ _01029_ _01028_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__o31a_1
X_15046_ _05940_ _05941_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__nand2_1
X_11209_ _02099_ _02119_ _02101_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__a21boi_2
XFILLER_96_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19854_ _00980_ _01069_ _01070_ VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__nand3_2
X_12189_ _03116_ _03119_ _03117_ net65 _03122_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__a311oi_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18805_ _09688_ _09692_ _09694_ VGND VGND VPWR VPWR _09698_ sky130_fd_sc_hd__a21o_1
X_16997_ _07863_ _07864_ _07865_ VGND VGND VPWR VPWR _07867_ sky130_fd_sc_hd__a21oi_1
X_19785_ _00888_ _00995_ _00889_ net407 VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__and4_1
X_15948_ net261 _06821_ _06823_ net262 VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__o211a_1
XFILLER_95_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18736_ net335 _09619_ _09598_ VGND VGND VPWR VPWR _09622_ sky130_fd_sc_hd__a21oi_1
XFILLER_48_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18667_ _09544_ _09546_ _09166_ _09329_ VGND VGND VPWR VPWR _09547_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15879_ net602 net527 VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__nand2_1
X_17618_ net1093 a_l\[11\] _02588_ VGND VGND VPWR VPWR _08482_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_65_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18598_ _09334_ _09462_ _09464_ _09466_ VGND VGND VPWR VPWR _09472_ sky130_fd_sc_hd__nand4_1
XFILLER_17_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17549_ _08411_ _08412_ _08293_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__and3_1
X_20560_ clknet_leaf_18_clk _00200_ VGND VGND VPWR VPWR mid_sum\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19219_ _10069_ _10114_ net206 _10008_ VGND VGND VPWR VPWR _10117_ sky130_fd_sc_hd__o211a_1
Xclkload9 clknet_leaf_60_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__bufinv_16
X_20491_ clknet_leaf_28_clk _00131_ VGND VGND VPWR VPWR term_mid\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ net646 net546 VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__nand2_1
X_20758_ clknet_leaf_52_clk _00398_ VGND VGND VPWR VPWR p_ll\[28\] sky130_fd_sc_hd__dfxtp_1
X_10511_ term_high\[56\] net1362 _01660_ _01662_ net796 VGND VGND VPWR VPWR _00073_
+ sky130_fd_sc_hd__a311oi_1
XFILLER_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11491_ _02428_ _02429_ _02336_ VGND VGND VPWR VPWR _02431_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13230_ net787 net784 net704 net700 VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__and4_1
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20689_ clknet_3_0__leaf_clk _00329_ VGND VGND VPWR VPWR p_hl\[23\] sky130_fd_sc_hd__dfxtp_2
X_10442_ net793 _01607_ _01608_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__and3_1
XFILLER_109_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13161_ _04080_ _04071_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nand2_1
X_10373_ _01311_ net444 _01439_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__a21oi_2
X_12112_ _03045_ _03046_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__nor2_1
X_13092_ _03958_ _03972_ _03973_ _04016_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__nand4_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16920_ _07788_ _07633_ _07787_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__nand3_2
X_12043_ net661 net508 VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__nand2_2
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16851_ _07446_ _07447_ _07444_ VGND VGND VPWR VPWR _07722_ sky130_fd_sc_hd__o21ai_2
X_15802_ net608 net601 VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__nand2_8
X_16782_ _07640_ _07647_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__nand2_1
X_19570_ _00758_ _00760_ net406 VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15733_ _06608_ _06599_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__nand2_1
X_18521_ _09364_ _09380_ _09382_ VGND VGND VPWR VPWR _09388_ sky130_fd_sc_hd__and3_1
XFILLER_46_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13994_ _09515_ _04897_ net656 _04896_ net778 VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__o2111ai_4
X_12945_ _03869_ _03870_ _03871_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__o21ai_1
X_15664_ _06540_ _06543_ _06541_ VGND VGND VPWR VPWR _06545_ sky130_fd_sc_hd__a21oi_2
X_18452_ _09305_ _09309_ _09205_ _09307_ VGND VGND VPWR VPWR _09313_ sky130_fd_sc_hd__o211a_4
X_12876_ net674 net474 _03799_ _03800_ VGND VGND VPWR VPWR _03804_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ net983 net706 net463 VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__and3_1
X_15595_ net616 net533 VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__nand2_1
X_17403_ _08163_ _08267_ _08268_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__nand3_2
X_18383_ net782 net1069 net573 net791 VGND VGND VPWR VPWR _09237_ sky130_fd_sc_hd__a22oi_4
X_14615_ _05514_ _05516_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__nand2_1
X_11758_ _02600_ _02602_ _02590_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a21oi_2
X_17334_ _08192_ _08194_ _08197_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_16_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _09220_ _09504_ _05271_ _05446_ _05445_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_60_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ p_hl\[13\] p_lh\[13\] VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__or2_1
X_11689_ net658 net525 net520 net664 VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__a22oi_4
X_17265_ _08083_ _08085_ _08131_ VGND VGND VPWR VPWR _08133_ sky130_fd_sc_hd__o21ai_1
X_19004_ _09890_ _09894_ VGND VGND VPWR VPWR _09895_ sky130_fd_sc_hd__nand2_2
X_14477_ b_l\[14\] net709 _05193_ _05191_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__a31o_1
X_16216_ _07002_ _07003_ _06994_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__o21a_1
X_17196_ _08051_ _08054_ _08057_ _07902_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a31oi_2
X_13428_ net766 net693 VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__nand2_1
X_16147_ _07020_ _07021_ _06953_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__nand3_4
XFILLER_114_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13359_ net763 net705 VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__nand2_1
XFILLER_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16078_ _06911_ _06912_ _06916_ _06893_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_75_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19906_ net574 net1043 net1099 net580 VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__a22o_1
X_15029_ net733 net657 VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_84_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19837_ _00895_ _01051_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__nand2_2
XFILLER_84_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 a[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19768_ _00975_ _00976_ _00970_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18719_ net887 net1082 VGND VGND VPWR VPWR _09604_ sky130_fd_sc_hd__nand2_1
X_19699_ net588 net729 net725 net591 VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__a22oi_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20612_ clknet_leaf_41_clk _00252_ VGND VGND VPWR VPWR p_ll_pipe\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20543_ clknet_leaf_44_clk _00183_ VGND VGND VPWR VPWR mid_sum\[6\] sky130_fd_sc_hd__dfxtp_1
X_20474_ clknet_leaf_42_clk _00114_ VGND VGND VPWR VPWR term_mid\[18\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_89_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_98_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10991_ _01906_ _01931_ _01932_ _01883_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_122_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ net321 _03656_ _03657_ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__nand3_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _03576_ _03578_ _03585_ _03586_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__nand4_1
X_11612_ _02471_ _02472_ _02546_ _02547_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _05126_ _05302_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__nand2_2
X_12592_ _03514_ _03520_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__nor2_1
XFILLER_51_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15380_ _06231_ _06227_ _06226_ _06225_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__a22o_1
XFILLER_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _09449_ _09602_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__nor2_1
Xwire400 _02365_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__buf_1
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14331_ _05050_ _05065_ _05223_ _05224_ _05063_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__o2111ai_2
XFILLER_128_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11474_ _02407_ _02408_ _02410_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__a21oi_1
XFILLER_109_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17050_ _07783_ net503 net1069 VGND VGND VPWR VPWR _07919_ sky130_fd_sc_hd__and3_1
X_14262_ _05158_ _05163_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__nand2_2
X_10425_ term_mid\[39\] term_high\[39\] _01592_ _01593_ VGND VGND VPWR VPWR _01594_
+ sky130_fd_sc_hd__a211o_1
X_16001_ net572 net542 VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__nand2_4
X_13213_ _04130_ _04132_ net65 VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__a21oi_1
X_14193_ _05095_ _05097_ _04960_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13144_ _04033_ _04038_ _04067_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__o21ai_1
X_10356_ term_low\[29\] term_mid\[29\] _01278_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__a21oi_1
X_17952_ _08803_ _08806_ _08800_ VGND VGND VPWR VPWR _08809_ sky130_fd_sc_hd__a21oi_1
X_10287_ _10148_ _10169_ _00482_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__nand3_1
X_13075_ _03904_ net885 net634 VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__and3_1
XFILLER_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12026_ _02960_ _02953_ _02809_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__o211a_1
X_16903_ _07766_ _07770_ _07772_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__a21o_1
X_17883_ _08742_ _08741_ VGND VGND VPWR VPWR _08743_ sky130_fd_sc_hd__nand2b_1
X_16834_ _07703_ _07704_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__nand2_1
Xclone323 net617 VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__clkbuf_16
X_19622_ _00606_ _00621_ _00608_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__o21ai_1
XFILLER_93_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16765_ _07633_ _07635_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__nor2_2
XFILLER_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19553_ net819 net562 net556 b_l\[6\] VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__a22oi_4
X_13977_ _04733_ _04875_ _04874_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a21o_1
X_16696_ _07450_ _07564_ _07565_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__nand3b_1
X_15716_ _06592_ _06594_ _06593_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__a21oi_4
XFILLER_74_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18504_ net780 net581 VGND VGND VPWR VPWR _09369_ sky130_fd_sc_hd__nand2_1
X_12928_ _03848_ _03851_ _03807_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__nand3_2
X_19484_ _00661_ _00662_ net408 VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__and3_1
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15647_ _06527_ _06523_ _06516_ _06526_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__o211ai_1
X_18435_ _09265_ _09266_ _09284_ _09287_ VGND VGND VPWR VPWR _09294_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_61_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12859_ _03782_ _03783_ _03712_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15578_ net797 _06457_ _06458_ _06459_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__nor4b_1
X_18366_ net1128 net1082 net737 net630 VGND VGND VPWR VPWR _09218_ sky130_fd_sc_hd__a22oi_1
XFILLER_147_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17317_ _02589_ _06867_ net600 net476 _08182_ VGND VGND VPWR VPWR _08184_ sky130_fd_sc_hd__o2111ai_4
X_18297_ net774 net769 net604 net1113 _09134_ VGND VGND VPWR VPWR _09143_ sky130_fd_sc_hd__a41o_1
X_14529_ _05303_ net670 net746 VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__and3_1
XFILLER_30_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17248_ _08112_ _08113_ net375 VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__nand3_4
Xmax_cap700 net701 VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__buf_12
X_17179_ _07812_ _07906_ _08045_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__a21oi_1
Xmax_cap722 net723 VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__clkbuf_8
Xmax_cap733 net736 VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__buf_8
Xmax_cap755 b_l\[7\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__buf_12
Xmax_cap766 net768 VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__buf_12
Xmax_cap788 net789 VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__buf_12
Xmax_cap777 net778 VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__buf_12
X_20190_ _01358_ _01378_ _01379_ _01427_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__nand4_2
XFILLER_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20526_ clknet_leaf_47_clk _00166_ VGND VGND VPWR VPWR term_low\[21\] sky130_fd_sc_hd__dfxtp_1
X_20457_ clknet_leaf_14_clk _00097_ VGND VGND VPWR VPWR term_high\[49\] sky130_fd_sc_hd__dfxtp_1
X_10210_ net957 VGND VGND VPWR VPWR _09471_ sky130_fd_sc_hd__clkinv_8
X_11190_ _02126_ _02128_ _02042_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_132_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20388_ clknet_leaf_41_clk _00028_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfxtp_1
XFILLER_88_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13900_ _04774_ _04776_ _04804_ _04805_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__o2bb2ai_2
X_14880_ _05658_ _05666_ _05778_ net65 VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__a31o_1
X_13831_ _04732_ _04734_ _04735_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__and3_1
X_16550_ net208 _07419_ _07309_ _07420_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__o211ai_2
X_10974_ _01918_ _01919_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__nand2_2
XFILLER_90_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13762_ net432 _04669_ _04668_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__o21ai_2
X_12713_ _09635_ _03639_ _03642_ VGND VGND VPWR VPWR _03643_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15501_ _06388_ _06389_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__xor2_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16481_ _07262_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__nand2_1
X_18220_ net781 net594 net585 net791 VGND VGND VPWR VPWR _09067_ sky130_fd_sc_hd__a22oi_2
XFILLER_70_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13693_ _04596_ _04597_ _04592_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a21o_1
X_12644_ _03534_ _03568_ _03569_ VGND VGND VPWR VPWR _03575_ sky130_fd_sc_hd__nand3_2
XFILLER_62_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15432_ _06323_ _06316_ _06322_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__nand3_1
X_18151_ _08997_ _08998_ _08963_ VGND VGND VPWR VPWR _08999_ sky130_fd_sc_hd__a21oi_2
X_12575_ _03432_ _03505_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__nand2_1
X_15363_ _06220_ _06253_ _06254_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__nand3_2
XFILLER_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11526_ _02463_ net712 _02461_ net483 VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__nand4_2
X_17102_ net451 _07970_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__nor2_1
X_18082_ _08910_ net374 _08928_ _08929_ VGND VGND VPWR VPWR _08931_ sky130_fd_sc_hd__o211ai_4
Xwire241 _06328_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__buf_1
Xwire230 _00548_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_6
XFILLER_8_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14314_ _05195_ _05197_ _05213_ _05215_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__a22o_1
X_17033_ net559 net554 net1023 net516 VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__and4_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire274 _00674_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__buf_1
X_15294_ _06122_ _06123_ _06090_ _06185_ _06186_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__a32o_1
XFILLER_144_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11457_ net686 net507 VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nand2_2
X_14245_ net767 net656 VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__nand2_1
X_10408_ term_mid\[38\] term_high\[38\] VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__and2_1
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11388_ _02131_ _02232_ _02140_ _02230_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__a31oi_1
X_14176_ _05072_ _05080_ _05079_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__o21ai_2
X_13127_ a_h\[13\] net641 net1150 net999 _04005_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__a41o_1
X_18984_ net621 net618 net729 net725 VGND VGND VPWR VPWR _09875_ sky130_fd_sc_hd__nand4_2
X_10339_ _01084_ _01095_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__or2_1
X_17935_ _08766_ _08768_ _08770_ _08777_ VGND VGND VPWR VPWR _08793_ sky130_fd_sc_hd__o22ai_1
X_13058_ _03981_ _03982_ _03977_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_55_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _02940_ net247 net712 net474 VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__o211ai_2
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17866_ _08629_ _08676_ _08686_ _08672_ _08682_ VGND VGND VPWR VPWR _08726_ sky130_fd_sc_hd__o221ai_4
XFILLER_39_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16817_ _07494_ _07499_ _07678_ _07681_ _07496_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__a221oi_1
XFILLER_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17797_ _08656_ _08646_ _08655_ VGND VGND VPWR VPWR _08659_ sky130_fd_sc_hd__nand3_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19605_ _00800_ _00801_ net588 net732 VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__nand4_2
X_16748_ _07597_ _07598_ _07614_ _07615_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__nand4_1
Xclone186 net1014 VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19536_ _09199_ _09384_ _00724_ _00725_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__o211ai_2
XFILLER_46_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _07546_ _07547_ _07509_ VGND VGND VPWR VPWR _07551_ sky130_fd_sc_hd__a21o_1
X_19467_ _00649_ _00650_ _00653_ _00455_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__o2bb2ai_2
X_18418_ net800 net610 net759 net754 VGND VGND VPWR VPWR _09276_ sky130_fd_sc_hd__nand4_1
X_19398_ _09188_ _09384_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__nor2_1
XFILLER_22_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18349_ _09087_ _09110_ _09198_ _09200_ VGND VGND VPWR VPWR _09201_ sky130_fd_sc_hd__a22oi_1
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20311_ _01555_ _01556_ net797 VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__a21oi_1
Xmax_cap530 b_h\[3\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_12
Xinput60 b[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20242_ _01484_ _01485_ _01457_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__and3b_1
Xmax_cap563 net564 VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__buf_12
Xmax_cap552 net553 VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__buf_8
XFILLER_143_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap596 a_l\[7\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__buf_8
XFILLER_103_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap585 net586 VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__buf_12
X_20173_ net727 net551 VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__nand2_1
Xmax_cap574 net576 VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__buf_12
XFILLER_131_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_97_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10690_ p_hl\[9\] p_lh\[9\] _01725_ _01726_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__o211ai_4
XFILLER_8_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ _03142_ _03143_ _03162_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_23_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11311_ _02155_ _02160_ _02157_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__a21o_1
XFILLER_5_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12291_ _03221_ _03222_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__nand2_1
X_20509_ clknet_leaf_32_clk _00149_ VGND VGND VPWR VPWR term_low\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_130_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11242_ _02182_ _02183_ _02153_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__a21oi_2
X_14030_ _04932_ _04933_ _04918_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__and3_1
XFILLER_134_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11173_ _02114_ _02115_ _02038_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__a21o_1
X_15981_ _06755_ _06767_ _06857_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__o21ai_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17720_ _08562_ _08575_ _08576_ _08377_ VGND VGND VPWR VPWR _08583_ sky130_fd_sc_hd__a31o_2
X_14932_ _05616_ _05716_ _05715_ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__o21a_1
XFILLER_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17651_ _08391_ _08406_ _08405_ VGND VGND VPWR VPWR _08515_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_50_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _05756_ _05758_ _05759_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__o21ai_1
X_16602_ _07471_ _07473_ net629 net477 VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__nand4b_2
XTAP_TAPCELL_ROW_50_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13814_ _04705_ _04714_ _04717_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__nand3_2
XFILLER_91_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17582_ _08429_ _08431_ _08439_ _08441_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__nand4_1
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14794_ _09493_ _09504_ _04260_ _09482_ _09264_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__o32a_1
X_19321_ net592 net738 VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__nand2_1
X_10957_ _01901_ _01865_ _01900_ _01880_ net796 VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__a41o_1
X_16533_ _07403_ _07404_ _07370_ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__a21oi_1
X_13745_ _04649_ net989 _04625_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__a21boi_2
X_16464_ _07318_ _07319_ _07330_ _07332_ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__o22ai_1
X_13676_ _04553_ _04565_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__nand2_2
X_19252_ _09994_ _10150_ _10149_ _10147_ VGND VGND VPWR VPWR _10153_ sky130_fd_sc_hd__o211ai_4
X_12627_ _03548_ _03549_ _03557_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a21oi_2
X_18203_ net769 net604 VGND VGND VPWR VPWR _09050_ sky130_fd_sc_hd__nand2_1
X_10888_ net794 net1256 VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__and2_1
X_15415_ _06304_ _06305_ _06301_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__a21oi_1
X_19183_ net609 net729 net725 net618 VGND VGND VPWR VPWR _10078_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16395_ _07110_ _07114_ _07111_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__a21oi_1
X_18134_ _08973_ _08974_ _08978_ VGND VGND VPWR VPWR _08982_ sky130_fd_sc_hd__nand3_2
X_12558_ _03357_ _03363_ VGND VGND VPWR VPWR _03490_ sky130_fd_sc_hd__nand2_1
X_15346_ _06238_ _06239_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__and2_1
X_11509_ _02424_ net269 _02423_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__a21boi_2
X_18065_ _08869_ _08872_ _08874_ VGND VGND VPWR VPWR _08914_ sky130_fd_sc_hd__o21ai_2
X_12489_ net1049 net633 b_h\[4\] net518 VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_57_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ _06159_ _06168_ _06170_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__and3_2
XFILLER_132_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17016_ _07863_ _07865_ _07864_ _07870_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__a31oi_1
X_14228_ _05125_ _05128_ net746 net676 VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__and4_1
XFILLER_125_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ net350 VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__inv_2
XFILLER_140_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18967_ _09856_ _09858_ VGND VGND VPWR VPWR _09859_ sky130_fd_sc_hd__nand2_1
X_17918_ _08773_ _08625_ _08775_ VGND VGND VPWR VPWR _08777_ sky130_fd_sc_hd__a21oi_4
X_18898_ _09680_ _09683_ _09685_ _09786_ _09787_ VGND VGND VPWR VPWR _09790_ sky130_fd_sc_hd__o2111ai_1
X_17849_ _08662_ _08707_ _08706_ VGND VGND VPWR VPWR _08710_ sky130_fd_sc_hd__a21o_1
XFILLER_82_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20791_ clknet_leaf_8_clk _00431_ VGND VGND VPWR VPWR a_l\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_81_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19519_ _10152_ _10153_ _00570_ _00571_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__and4_1
XFILLER_35_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer204 net753 VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__buf_4
XFILLER_147_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer237 _02907_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer215 net1009 VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_20_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer248 net617 VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__buf_6
Xrebuffer259 _05178_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap360 _02301_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_1
Xmax_cap371 _09240_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_1
XFILLER_1_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20225_ _01466_ _01467_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__nand2_1
XFILLER_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap393 _04641_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_4
XFILLER_89_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20156_ _01321_ _01332_ _01391_ _01394_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_76_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20087_ _01201_ _01246_ _01248_ _01319_ _01320_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__a32o_2
XFILLER_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11860_ _02761_ _02796_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__nand2_1
XFILLER_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ net664 net518 _02724_ _02726_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__a22o_1
X_10811_ p_hl\[28\] p_lh\[28\] VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__and2_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _01768_ _01770_ _01765_ _01766_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__a211oi_1
X_13530_ net751 net705 VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__nand2_1
XFILLER_26_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10673_ _01712_ _01710_ _01709_ net797 VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__a31o_1
X_13461_ _04371_ _04319_ _04370_ VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__nand3_2
XFILLER_9_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15200_ net739 net733 net909 a_h\[14\] VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__nand4_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16180_ _07055_ _07054_ net797 VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__a21oi_1
X_12412_ _03169_ _03209_ _03211_ _03170_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__a31oi_4
X_13392_ _04268_ _04302_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__nand3b_4
XFILLER_138_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12343_ _03268_ _03269_ _03254_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__a21o_1
X_15131_ _06019_ _06020_ _06018_ VGND VGND VPWR VPWR _06028_ sky130_fd_sc_hd__o21a_1
XFILLER_126_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12274_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03208_ sky130_fd_sc_hd__a21o_1
X_15062_ _05920_ _05955_ _05957_ VGND VGND VPWR VPWR _05960_ sky130_fd_sc_hd__nand3_2
X_11225_ net664 net965 VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__nand2_1
X_14013_ _04734_ _04735_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__nand2_1
XFILLER_134_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19870_ _01065_ _01055_ _01054_ VGND VGND VPWR VPWR _01087_ sky130_fd_sc_hd__o21a_1
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ _02098_ _02061_ _02097_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__nand3_2
XFILLER_110_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18821_ _09530_ _09562_ _09528_ VGND VGND VPWR VPWR _09714_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_52_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11087_ _02026_ _02027_ _02015_ _02017_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__o211ai_1
XFILLER_110_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15964_ net173 _06836_ _06839_ _06840_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__o211ai_4
X_18752_ net775 net576 VGND VGND VPWR VPWR _09640_ sky130_fd_sc_hd__nand2_1
X_17703_ net550 net500 net494 net555 VGND VGND VPWR VPWR _08566_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14915_ _05806_ _05808_ _05810_ VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__and3_1
X_15895_ net583 net1063 net521 net607 VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__a22oi_1
XFILLER_76_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18683_ _09529_ _09530_ _09562_ VGND VGND VPWR VPWR _09565_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17634_ _08395_ _08494_ net565 net488 _08493_ VGND VGND VPWR VPWR _08498_ sky130_fd_sc_hd__o2111ai_4
X_14846_ _05708_ _05741_ _05743_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__nand3_2
XFILLER_17_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17565_ _08299_ _08374_ _08426_ _08428_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_67_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14777_ _05675_ _05676_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__nor2_1
X_11989_ _02924_ _02860_ _02923_ VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__nand3_4
X_16516_ _07381_ _07382_ _07386_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__nand3_2
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13728_ net757 net752 net694 net689 VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__and4_1
XFILLER_16_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19304_ net1065 _00469_ _00470_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__and3_1
X_17496_ _08248_ _08253_ _08360_ _08359_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__a22o_1
X_19235_ _10132_ _10120_ VGND VGND VPWR VPWR _10134_ sky130_fd_sc_hd__nand2_1
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16447_ _07318_ _07319_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ _04551_ _04553_ net288 VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand3_2
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16378_ _07247_ _07250_ _07240_ _07241_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__o211ai_1
X_19166_ _10057_ _10033_ _10056_ _09938_ VGND VGND VPWR VPWR _10059_ sky130_fd_sc_hd__nand4_4
X_18117_ net779 net605 VGND VGND VPWR VPWR _08965_ sky130_fd_sc_hd__nand2_1
X_19097_ _09976_ _09977_ _09987_ VGND VGND VPWR VPWR _09988_ sky130_fd_sc_hd__a21o_4
XFILLER_8_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15329_ _06221_ _06222_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__nand2_1
X_18048_ net805 _06441_ _08863_ _08895_ VGND VGND VPWR VPWR _08897_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_6_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20010_ _01232_ _01233_ _01215_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__a21o_1
XFILLER_101_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19999_ _01224_ _01216_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__nand2_1
XFILLER_104_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_61_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20774_ clknet_leaf_0_clk _00414_ VGND VGND VPWR VPWR a_h\[12\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_98_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 mid_sum\[27\] VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold471 p_ll\[12\] VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold482 p_hh_pipe\[22\] VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 p_hh_pipe\[20\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _01950_ _01951_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__nand2_1
XFILLER_104_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20208_ _01443_ _01446_ _01449_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_129_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20139_ _09351_ _01370_ net721 net568 _01372_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__o2111ai_4
XTAP_TAPCELL_ROW_142_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12961_ _09471_ _09679_ _03881_ _03882_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__o211a_1
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11912_ _02843_ _02845_ net399 VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__a21o_1
X_15680_ _06493_ _06433_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__nand2_1
X_12892_ _03744_ _03749_ _03747_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__a21o_1
X_14700_ _05432_ _05428_ _05424_ _05429_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__o2bb2ai_4
X_11843_ _02777_ _02769_ _02776_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__nand3_2
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14631_ _05530_ _05528_ _05405_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_107_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _08215_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__nand2_1
XFILLER_14_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16301_ _07045_ _07173_ _07170_ net161 VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__o211a_1
X_11774_ _02650_ _02707_ net682 net501 _02706_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__o2111ai_2
X_14562_ _05460_ _05415_ _05459_ _05297_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__nand4_4
XPHY_EDGE_ROW_109_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17281_ _07892_ net419 _07890_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__a21oi_4
X_10725_ p_hl\[15\] p_lh\[15\] p_hl\[14\] p_lh\[14\] VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__o211a_1
X_13513_ _04349_ _04416_ net777 net675 _04415_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o2111ai_1
X_14493_ _05377_ _05391_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__nand2_1
X_16232_ _06982_ _07092_ _07103_ _07105_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__o22a_1
X_10656_ p_hl\[5\] p_lh\[5\] VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__nand2_1
X_13444_ _04351_ _04352_ _04348_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__a21o_1
X_19020_ net760 net753 net589 net580 VGND VGND VPWR VPWR _09911_ sky130_fd_sc_hd__nand4_1
X_16163_ _06954_ _07018_ _07019_ net259 VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__a31oi_2
Xclkload16 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__inv_12
Xclkload38 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__inv_12
X_10587_ net793 net1222 VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__and2_1
Xclkload49 clknet_leaf_39_clk VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__inv_12
X_13375_ net784 net675 VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15114_ net726 net723 net958 net663 VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__nand4_1
Xclkload27 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_16
X_16094_ _09144_ _09613_ _06794_ _06901_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__o22a_1
XFILLER_126_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12326_ net647 net511 net508 net906 VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__a22oi_1
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12257_ _03186_ _03187_ net682 net489 VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__nand4_1
XFILLER_79_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19922_ _01009_ _01011_ _01029_ _01028_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__o31ai_1
X_15045_ net726 net723 net862 net668 VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__nand4_2
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12188_ _03119_ _03117_ _03116_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__and3_1
X_11208_ _02099_ _02119_ _02100_ _02095_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_79_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19853_ _01057_ _01065_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18804_ _09688_ _09692_ _09694_ VGND VGND VPWR VPWR _09697_ sky130_fd_sc_hd__a21oi_1
X_16996_ _07704_ _07712_ _07703_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__a21boi_1
X_11139_ net678 net671 VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__nand2_8
X_19784_ _00992_ net366 _00991_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__a21oi_2
X_15947_ _06823_ net262 VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__nand2_1
X_18735_ _09614_ _09618_ _09598_ net925 VGND VGND VPWR VPWR _09621_ sky130_fd_sc_hd__o211ai_4
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15878_ net587 net541 VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__nand2_1
XFILLER_64_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18666_ _09540_ _09541_ _09531_ VGND VGND VPWR VPWR _09546_ sky130_fd_sc_hd__nand3_2
X_17617_ a_l\[11\] net485 VGND VGND VPWR VPWR _08481_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14829_ _05726_ _05727_ _05714_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__a21o_1
XFILLER_36_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18597_ _09462_ _09464_ _09465_ _09333_ VGND VGND VPWR VPWR _09470_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_127_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17548_ _08294_ _08409_ _08410_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__nand3_2
X_17479_ _08115_ _08119_ _08195_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__o21ai_1
X_20490_ clknet_leaf_18_clk _00130_ VGND VGND VPWR VPWR term_mid\[34\] sky130_fd_sc_hd__dfxtp_1
X_19218_ _10070_ _10071_ _10110_ _10112_ VGND VGND VPWR VPWR _10116_ sky130_fd_sc_hd__nand4_1
XFILLER_118_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19149_ net765 net567 VGND VGND VPWR VPWR _10041_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_584 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_145_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20757_ clknet_leaf_52_clk _00397_ VGND VGND VPWR VPWR p_ll\[27\] sky130_fd_sc_hd__dfxtp_1
X_10510_ term_high\[56\] _01660_ net1362 VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__a21oi_1
X_11490_ _02429_ _02336_ _02428_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__nand3_2
X_10441_ _01606_ _01603_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__nand2_1
XFILLER_108_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire626 net627 VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__buf_12
Xwire648 a_h\[12\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__buf_12
XFILLER_11_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20688_ clknet_3_0__leaf_clk _00328_ VGND VGND VPWR VPWR p_hl\[22\] sky130_fd_sc_hd__dfxtp_2
XFILLER_136_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13160_ _04080_ _04082_ _04071_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__a21o_1
X_10372_ _01311_ _01450_ _01428_ _01364_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__a211o_4
XFILLER_123_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12111_ net706 net475 _03042_ _03044_ VGND VGND VPWR VPWR _03046_ sky130_fd_sc_hd__a22oi_4
X_13091_ _03891_ _03959_ _03963_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_123_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12042_ _02864_ _02976_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__nand2_1
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16850_ _07718_ _07720_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__nand2_1
XFILLER_49_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15801_ _06678_ _06679_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__nand2_2
X_16781_ _07641_ _07642_ _07640_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__o21a_2
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13993_ _09515_ _04897_ _04891_ _04896_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__o211a_1
X_15732_ _09231_ _09581_ net1070 _06605_ _06604_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__o221ai_4
X_12944_ _03869_ _03870_ _03782_ _03784_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__o211a_1
X_18520_ _09386_ VGND VGND VPWR VPWR _09387_ sky130_fd_sc_hd__inv_2
XFILLER_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18451_ net1042 _09310_ _09311_ VGND VGND VPWR VPWR _09312_ sky130_fd_sc_hd__nand3_2
XFILLER_34_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15663_ _06536_ _06537_ _06543_ VGND VGND VPWR VPWR _06544_ sky130_fd_sc_hd__o21ai_1
X_17402_ _08267_ _08268_ _08163_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__a21o_1
X_12875_ _03799_ _03800_ _03801_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__a21o_1
XFILLER_65_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11826_ net706 net483 net481 net708 VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__a22o_1
X_15594_ net625 net528 VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__nand2_1
X_18382_ net791 net573 VGND VGND VPWR VPWR _09236_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _05510_ _05512_ _05509_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__a21o_1
X_11757_ _02598_ _02601_ _02600_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__o21a_1
X_17333_ _08193_ _08195_ _08197_ VGND VGND VPWR VPWR _08200_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_16_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _05442_ _05443_ _05446_ _05271_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__o2bb2ai_1
X_17264_ _08127_ net235 _08084_ _08086_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_60_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ p_hl\[13\] p_lh\[13\] VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__nand2_1
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16215_ _06974_ _07014_ _07015_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__a21oi_1
X_11688_ net672 net518 VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__nand2_1
X_19003_ _09891_ _09884_ _09881_ _09892_ VGND VGND VPWR VPWR _09894_ sky130_fd_sc_hd__o211ai_2
X_14476_ b_l\[15\] net709 VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__nand2_1
X_10639_ _01676_ _01678_ _01683_ net797 VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__a31o_1
X_17195_ _08059_ _07902_ _08058_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__nand3_4
X_13427_ net772 net766 net693 net986 VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand4_4
XFILLER_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16146_ _06893_ _06918_ _07018_ _07019_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__o211ai_4
X_13358_ _04241_ _04232_ _04230_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__a21oi_1
X_16077_ _06894_ _06913_ _06915_ _06890_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__o2bb2ai_2
X_12309_ _03238_ _03240_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__nand2_1
XFILLER_114_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13289_ _04189_ _04200_ _04201_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__nand3_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19905_ net589 net721 VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__nand2_1
X_15028_ net739 net651 VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__nand2_1
XFILLER_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19836_ _00943_ _00938_ _00894_ _00945_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__o211ai_2
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19767_ _10005_ _00712_ _00973_ _00976_ _00970_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__o311a_1
X_16979_ _07844_ _07842_ _07734_ _07697_ _07847_ VGND VGND VPWR VPWR _07849_ sky130_fd_sc_hd__a221oi_2
Xinput3 a[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_18718_ net619 net737 VGND VGND VPWR VPWR _09603_ sky130_fd_sc_hd__nand2_1
X_19698_ net591 net588 net729 net725 VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__nand4_2
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18649_ _09524_ _09525_ _09445_ VGND VGND VPWR VPWR _09528_ sky130_fd_sc_hd__a21oi_1
XFILLER_25_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20611_ clknet_leaf_36_clk _00251_ VGND VGND VPWR VPWR p_ll_pipe\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20542_ clknet_leaf_43_clk _00182_ VGND VGND VPWR VPWR mid_sum\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20473_ clknet_leaf_37_clk _00113_ VGND VGND VPWR VPWR term_mid\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10990_ _01932_ _01906_ _01931_ _01883_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_122_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _03576_ _03578_ _03587_ VGND VGND VPWR VPWR _03591_ sky130_fd_sc_hd__nand3_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _02475_ _02547_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__nand2_1
X_20809_ clknet_leaf_0_clk _00449_ VGND VGND VPWR VPWR b_h\[15\] sky130_fd_sc_hd__dfxtp_4
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ net353 _03516_ _03519_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_13_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _05223_ _05224_ _05226_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_137_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire401 _02346_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_1
XFILLER_128_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11542_ _02367_ _02371_ _02382_ _02369_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__o22ai_2
Xwire423 _06436_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_1
Xwire412 _09652_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ _02407_ _02408_ _02409_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__nand3_1
Xwire434 _04347_ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14261_ _05163_ net643 net778 VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__nand3_1
X_10424_ term_mid\[39\] term_high\[39\] term_mid\[38\] term_high\[38\] VGND VGND VPWR
+ VPWR _01593_ sky130_fd_sc_hd__o211a_1
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16000_ net966 net521 VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__nand2_1
X_13212_ _04097_ _04098_ _04117_ _04119_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__o22a_1
X_14192_ _04953_ _04957_ _05093_ _05094_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__a22o_1
XFILLER_109_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ _04065_ _04066_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10355_ term_low\[29\] term_mid\[29\] term_low\[28\] term_mid\[28\] VGND VGND VPWR
+ VPWR _01278_ sky130_fd_sc_hd__o211a_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17951_ _08776_ _08804_ _08802_ net170 VGND VGND VPWR VPWR _08808_ sky130_fd_sc_hd__a211oi_1
X_13074_ _03997_ _03998_ _03999_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__o21a_1
X_10286_ term_low\[20\] term_mid\[20\] VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__nand2_1
XFILLER_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12025_ _02956_ _02695_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__nand2_1
X_16902_ _07600_ _07610_ _07611_ _07599_ _07614_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__a32o_2
XFILLER_104_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17882_ _08701_ _08703_ _08702_ VGND VGND VPWR VPWR _08742_ sky130_fd_sc_hd__a21boi_1
X_16833_ _07591_ _07702_ _07701_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__nand3_2
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19621_ _00617_ _00618_ _00607_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__o21a_1
X_16764_ net566 net523 net516 net571 VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__a22oi_2
XFILLER_80_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19552_ net1121 net755 net562 net556 VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__nand4_4
X_13976_ _04733_ _04875_ _04874_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__a21oi_1
X_16695_ _07566_ _07450_ VGND VGND VPWR VPWR _07567_ sky130_fd_sc_hd__nand2_1
X_15715_ _06592_ _06591_ net624 net515 VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__and4_1
XFILLER_73_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18503_ _09234_ _09239_ _09237_ VGND VGND VPWR VPWR _09368_ sky130_fd_sc_hd__a21oi_1
X_12927_ _09613_ _03806_ _03853_ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__o211ai_2
X_19483_ _00661_ net833 net408 VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__a21o_1
X_15646_ _06440_ _06521_ _06518_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__o21ai_2
X_12858_ _03712_ _03782_ _03783_ VGND VGND VPWR VPWR _03787_ sky130_fd_sc_hd__nand3_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18434_ _09265_ _09266_ _09285_ _09288_ VGND VGND VPWR VPWR _09293_ sky130_fd_sc_hd__nand4_1
X_11809_ _02742_ _02743_ _02731_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__nand3_4
X_18365_ net1128 net630 net1082 VGND VGND VPWR VPWR _09217_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_32_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15577_ _06425_ _06454_ _06455_ _06410_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__and4_1
X_17316_ _02589_ _06867_ net600 net476 _08182_ VGND VGND VPWR VPWR _08183_ sky130_fd_sc_hd__o2111a_1
X_12789_ _03627_ _03630_ _03661_ _03667_ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__o22a_1
XFILLER_147_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18296_ _09136_ _09138_ _09199_ _09220_ VGND VGND VPWR VPWR _09142_ sky130_fd_sc_hd__o2bb2ai_1
X_14528_ _05417_ _05423_ _05425_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__nand3_1
X_17247_ _08114_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__inv_2
X_14459_ _05360_ _05137_ _05359_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__nand3_4
XFILLER_134_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap712 net713 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__buf_8
XFILLER_127_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17178_ _09373_ _09592_ _07645_ _07906_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_77_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16129_ _09231_ _09602_ _06589_ _06999_ _06998_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__o221a_1
Xmax_cap723 b_l\[13\] VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__buf_8
Xmax_cap745 net746 VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__buf_12
Xmax_cap734 net735 VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__buf_12
XFILLER_103_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap756 net758 VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__buf_12
Xmax_cap767 net768 VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19819_ _01009_ _01011_ _01028_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__o21ai_2
XFILLER_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_30 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20525_ clknet_leaf_43_clk _00165_ VGND VGND VPWR VPWR term_low\[20\] sky130_fd_sc_hd__dfxtp_1
X_20456_ clknet_leaf_15_clk _00096_ VGND VGND VPWR VPWR term_high\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_115_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20387_ clknet_leaf_41_clk _00027_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13830_ _04732_ _04734_ net762 net676 VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__and4_1
X_10973_ net686 net545 VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__nand2_2
XFILLER_56_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13761_ _04661_ _04663_ _04664_ _04556_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__a31o_1
XFILLER_16_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16480_ net590 net513 VGND VGND VPWR VPWR _07353_ sky130_fd_sc_hd__nand2_2
X_12712_ _03637_ _03638_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__nand2_1
XFILLER_71_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15500_ _06368_ _06374_ _06376_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13692_ _09155_ _09471_ _02362_ _04134_ _04596_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__o221ai_2
X_15431_ net716 net650 _06320_ _06321_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__a22o_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12643_ _03568_ _03569_ _03534_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__a21o_1
XFILLER_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18150_ _08992_ _08993_ _08980_ _08982_ VGND VGND VPWR VPWR _08998_ sky130_fd_sc_hd__o211ai_4
X_12574_ net638 net514 VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__nand2_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15362_ _06220_ _06253_ _06254_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__and3_1
X_11525_ _02461_ _02463_ _09177_ _09657_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__o2bb2ai_2
X_17101_ net606 net600 net485 net479 _07966_ VGND VGND VPWR VPWR _07970_ sky130_fd_sc_hd__a41o_1
X_18081_ _08928_ _08929_ VGND VGND VPWR VPWR _08930_ sky130_fd_sc_hd__nand2_1
Xwire231 _09636_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_1
XFILLER_8_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14313_ _05195_ _05197_ _05213_ _05215_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__nand4_2
X_15293_ _06122_ _06123_ _06090_ _06185_ _06186_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__a32oi_4
X_17032_ net554 net523 net516 net558 VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__a22o_1
X_14244_ net771 net650 VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__nand2_1
XFILLER_137_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11456_ _02255_ _02395_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_59_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire286 _04672_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__buf_1
Xwire297 _00592_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
X_10407_ term_mid\[38\] term_high\[38\] VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__nor2_1
X_11387_ net200 _02325_ net179 VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o21ai_2
X_14175_ _05068_ _05069_ _05040_ net316 VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__a31o_1
X_13126_ _09515_ _09657_ _04002_ _04006_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__o31a_1
X_18983_ net621 net618 _05043_ VGND VGND VPWR VPWR _09874_ sky130_fd_sc_hd__and3_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10338_ term_low\[28\] term_mid\[28\] VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__and2_1
XFILLER_124_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17934_ _08791_ VGND VGND VPWR VPWR _08792_ sky130_fd_sc_hd__inv_2
XFILLER_79_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _03981_ _03982_ net1019 b_h\[15\] VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__nand4_2
X_12008_ _02940_ net247 net712 net474 VGND VGND VPWR VPWR _02944_ sky130_fd_sc_hd__o211a_1
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10269_ _10018_ _10072_ VGND VGND VPWR VPWR _10083_ sky130_fd_sc_hd__or2_1
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17865_ net961 net555 net486 net999 _08681_ VGND VGND VPWR VPWR _08725_ sky130_fd_sc_hd__a41o_1
X_16816_ _07678_ _07681_ _07683_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__and3_1
X_17796_ _08647_ _08654_ _08646_ VGND VGND VPWR VPWR _08658_ sky130_fd_sc_hd__a21boi_1
X_19604_ net588 net732 VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__nand2_1
X_16747_ _07597_ _07598_ _07614_ _07615_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__a22o_1
XFILLER_93_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclone198 net1022 VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__clkbuf_16
XFILLER_81_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19535_ _09199_ _09384_ _00724_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__o21ai_2
XFILLER_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13959_ _04863_ _04864_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__nand2_1
XFILLER_81_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16678_ _07549_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__inv_2
X_19466_ net755 net562 VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__nand2_4
X_15629_ _06507_ _06509_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__nand2_1
X_18417_ _09271_ _09272_ VGND VGND VPWR VPWR _09274_ sky130_fd_sc_hd__nand2_2
X_19397_ _00554_ _00542_ _00544_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__a21boi_4
X_18348_ _09182_ _09185_ _09191_ _09193_ VGND VGND VPWR VPWR _09200_ sky130_fd_sc_hd__nand4_2
X_18279_ _09122_ _09123_ _09114_ VGND VGND VPWR VPWR _09125_ sky130_fd_sc_hd__a21o_1
XFILLER_147_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20310_ net1102 b_l\[14\] net548 b_l\[15\] _01546_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__a41oi_1
Xinput50 b[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 b[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xmax_cap542 net543 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__buf_12
Xmax_cap531 net533 VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__buf_12
X_20241_ _01484_ _01485_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__and2b_1
XFILLER_131_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap586 net587 VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__buf_12
XFILLER_107_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap597 net599 VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__buf_12
Xmax_cap564 net565 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__buf_12
Xmax_cap575 net576 VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__buf_8
X_20172_ net557 net724 VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__nand2_1
XFILLER_115_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11310_ _02186_ _02212_ _02184_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__a21oi_4
XFILLER_21_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12290_ _03068_ _03078_ _03221_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__and3_1
X_20508_ clknet_leaf_33_clk _00148_ VGND VGND VPWR VPWR term_low\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_113_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20439_ clknet_leaf_13_clk _00079_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11241_ net1046 _02162_ _02176_ _02177_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__o211ai_4
X_11172_ _02111_ _02105_ _02103_ _02110_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__o211ai_4
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15980_ _06776_ _06777_ _06769_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__o21ai_1
XFILLER_121_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14931_ _09308_ _09471_ _05824_ _05825_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_145_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17650_ _08391_ _08405_ VGND VGND VPWR VPWR _08514_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_50_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14862_ _05756_ _05758_ _05759_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__o21a_1
X_16601_ net840 net620 net484 net480 VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__nand4_2
X_17581_ _08429_ _08431_ _08442_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__a21o_1
X_13813_ _04704_ _04714_ _04717_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16532_ _07241_ _07368_ _07402_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__nand3_1
X_14793_ _05679_ _05686_ _05687_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__nand3_2
X_19320_ net598 net732 VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__nand2_1
X_10956_ _01882_ _01902_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__or2_1
X_13744_ net989 _04649_ _04619_ _04624_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_43_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16463_ _07320_ _07331_ _07333_ VGND VGND VPWR VPWR _07336_ sky130_fd_sc_hd__nand3_1
X_13675_ _09690_ _04582_ _04583_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__and3_1
X_10887_ net794 net1247 VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__and2_1
X_19251_ _10145_ _10146_ _10151_ VGND VGND VPWR VPWR _10152_ sky130_fd_sc_hd__nand3_1
XFILLER_31_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16394_ net950 net515 _06694_ _07113_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__o2bb2a_1
X_12626_ _03555_ _03556_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__nand2_1
X_18202_ net610 net769 net605 net774 VGND VGND VPWR VPWR _09049_ sky130_fd_sc_hd__a22oi_4
X_15414_ _06301_ _06304_ _06305_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__and3_1
X_19182_ net618 net609 net729 net725 VGND VGND VPWR VPWR _10077_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_42_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18133_ _08974_ _08978_ VGND VGND VPWR VPWR _08981_ sky130_fd_sc_hd__nand2_1
X_15345_ _06157_ _06175_ _06235_ _06236_ _06172_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12557_ _03485_ net176 _03376_ _03484_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__o211ai_4
XFILLER_8_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11508_ _02423_ _02427_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__nand2_1
X_18064_ _08910_ _08912_ VGND VGND VPWR VPWR _08913_ sky130_fd_sc_hd__nor2_4
X_12488_ net633 net518 VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__nand2_1
X_15276_ _06159_ _06170_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__nand2_1
X_17015_ _07882_ _07883_ _07884_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__o21a_1
X_11439_ net681 net517 _02376_ _02377_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__a22o_1
X_14227_ net746 net676 _05125_ _05128_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__a22o_1
XFILLER_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14158_ _04843_ _04851_ _05061_ _05062_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__o211ai_4
XFILLER_140_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13109_ _03949_ _03997_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__nand2_1
XFILLER_140_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18966_ _09716_ _09722_ _09854_ _09855_ VGND VGND VPWR VPWR _09858_ sky130_fd_sc_hd__a22o_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14089_ _04981_ _04991_ _04992_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nand3_1
X_17917_ _08774_ _08624_ _08775_ VGND VGND VPWR VPWR _08776_ sky130_fd_sc_hd__o21bai_2
XFILLER_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18897_ _09786_ _09787_ _09788_ VGND VGND VPWR VPWR _09789_ sky130_fd_sc_hd__a21bo_1
X_17848_ _08708_ VGND VGND VPWR VPWR _08709_ sky130_fd_sc_hd__inv_2
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17779_ _08632_ _08633_ _08638_ _08640_ VGND VGND VPWR VPWR _08641_ sky130_fd_sc_hd__a22o_1
XFILLER_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20790_ clknet_leaf_8_clk _00430_ VGND VGND VPWR VPWR a_l\[12\] sky130_fd_sc_hd__dfxtp_4
X_19518_ _00707_ _00708_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__nand2_1
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19449_ _00629_ _00632_ _00631_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__o21ai_1
Xrebuffer205 _00682_ VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__buf_1
Xrebuffer238 _02928_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer227 net536 VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlymetal6s4s_1
XTAP_TAPCELL_ROW_20_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer249 _02161_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__buf_2
XFILLER_147_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap361 _02200_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_112_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap372 _09071_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_4
XFILLER_2_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20224_ _01465_ _01458_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__or2_1
Xmax_cap350 _05063_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_2
Xmax_cap383 net384 VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap394 _03962_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
X_20155_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__inv_2
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20086_ _01234_ net330 _01309_ _01314_ _01316_ VGND VGND VPWR VPWR _01320_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_127_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ net665 net518 VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__nand2_1
X_10810_ p_hl\[28\] p_lh\[28\] VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__nor2_1
XFILLER_41_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ _01768_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__nand2_1
XFILLER_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13460_ _04365_ _04366_ _04333_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a21o_1
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12411_ _03295_ _03298_ _03336_ _03340_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__o2bb2ai_1
X_10672_ _01709_ _01710_ _01712_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_20_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_13391_ _04269_ _04297_ _04298_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__nand3_2
XFILLER_139_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12342_ _03268_ _03269_ _03253_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__nand3_2
X_15130_ _06021_ _06023_ _06018_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__a21o_1
XFILLER_126_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12273_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__a21oi_1
X_15061_ _05957_ _05919_ VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__nand2_2
XFILLER_135_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11224_ net671 net539 VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__nand2_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14012_ net746 _04711_ net694 _04709_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_147_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11155_ _02091_ _02092_ _02073_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__a21o_1
X_18820_ _09630_ _09631_ _09707_ _09708_ VGND VGND VPWR VPWR _09713_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15963_ _06728_ _06832_ _06835_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__and3_1
X_11086_ net403 _02025_ _02015_ _02017_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__o211ai_2
XFILLER_67_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18751_ net763 net942 VGND VGND VPWR VPWR _09639_ sky130_fd_sc_hd__nand2_1
X_17702_ net550 net500 VGND VGND VPWR VPWR _08565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14914_ _05806_ _05808_ _05809_ VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__nand3_2
X_15894_ net583 net1063 VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__nand2_1
XFILLER_64_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18682_ _09529_ _09530_ _09558_ _09561_ VGND VGND VPWR VPWR _09564_ sky130_fd_sc_hd__nand4_2
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17633_ net565 net488 VGND VGND VPWR VPWR _08497_ sky130_fd_sc_hd__nand2_1
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14845_ _05706_ _05707_ _05741_ _05743_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__nand4_4
X_11988_ _02877_ _02879_ _02916_ _02917_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__a22o_1
X_17564_ _08299_ _08374_ _08426_ _08428_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_67_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14776_ net761 net640 net636 net767 VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__a22oi_1
X_10939_ net697 net538 VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__nand2_1
X_16515_ _07372_ _07379_ _07386_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__o21ai_1
XFILLER_16_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19303_ net1065 _00469_ _00470_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__a21o_1
X_13727_ net752 net689 VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__nand2_2
X_17495_ _08252_ _08249_ _08247_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__o21ai_1
X_19234_ _10129_ _10131_ VGND VGND VPWR VPWR _10133_ sky130_fd_sc_hd__nand2_1
X_16446_ _07313_ _07315_ a_l\[0\] net477 VGND VGND VPWR VPWR _07319_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_80_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13658_ _04551_ net288 VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__nand2_4
X_16377_ _07242_ _07249_ _07248_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_11_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12609_ net1015 net995 net495 net659 VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__a22oi_1
X_13589_ _04492_ _04495_ _04496_ _04405_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__o2bb2ai_2
X_19165_ _10055_ _09951_ _10054_ _09937_ VGND VGND VPWR VPWR _10058_ sky130_fd_sc_hd__nand4_4
X_18116_ _08913_ _08929_ _08928_ VGND VGND VPWR VPWR _08964_ sky130_fd_sc_hd__a21boi_1
X_19096_ _09984_ _09986_ VGND VGND VPWR VPWR _09987_ sky130_fd_sc_hd__nand2_1
X_15328_ net722 net650 VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__nand2_1
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18047_ net922 _06441_ _08858_ _08862_ VGND VGND VPWR VPWR _08896_ sky130_fd_sc_hd__o22a_4
X_15259_ net719 net1019 _06150_ _06152_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__a22o_1
XFILLER_133_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19998_ _09308_ _09319_ _01110_ _01218_ _01223_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__o221ai_4
X_18949_ _09791_ _09792_ _09835_ _09837_ VGND VGND VPWR VPWR _09841_ sky130_fd_sc_hd__nand4_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20773_ clknet_leaf_0_clk _00413_ VGND VGND VPWR VPWR a_h\[11\] sky130_fd_sc_hd__dfxtp_4
XFILLER_136_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold461 p_hh_pipe\[15\] VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 p_hh_pipe\[23\] VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap180 _02138_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__buf_6
XFILLER_104_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold450 p_ll\[15\] VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 p_hh\[18\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold494 p_hh\[23\] VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap191 _06635_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_2
X_20207_ _01396_ _01398_ _01445_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_129_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20138_ _09351_ _01370_ _01368_ _01372_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__o211a_1
X_12960_ _03881_ _03882_ _03879_ VGND VGND VPWR VPWR _03887_ sky130_fd_sc_hd__a21o_1
XFILLER_58_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20069_ _01221_ _01294_ net731 net557 _01298_ VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_142_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ net399 _02843_ _02845_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__nand3_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12891_ _03815_ _03817_ VGND VGND VPWR VPWR _03819_ sky130_fd_sc_hd__nand2_1
X_11842_ _02773_ _02775_ _02770_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__a21o_1
XFILLER_73_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14630_ _05395_ _05404_ _05527_ _05529_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_107_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _05462_ _05322_ _05461_ _05298_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__nand4_4
X_16300_ _07174_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__inv_2
X_11773_ _02706_ _02709_ _09439_ _09613_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__o2bb2ai_1
X_13512_ net433 _04419_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nand2_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17280_ _08145_ _08147_ VGND VGND VPWR VPWR _08148_ sky130_fd_sc_hd__nand2_1
X_10724_ p_hl\[13\] p_lh\[13\] _01755_ _01748_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__o211ai_4
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14492_ _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__inv_2
X_16231_ _09592_ _07101_ net540 _07099_ net570 VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__o2111ai_2
X_10655_ _01691_ _01694_ _01693_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13443_ net787 net785 net675 net673 _04348_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__a41o_1
XFILLER_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16162_ _07025_ _07037_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__nand2_1
XFILLER_139_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13374_ _04221_ _04284_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__nand2_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload17 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__inv_16
Xclkload39 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__inv_8
X_10586_ net793 net1231 VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__and2_1
Xclkload28 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__clkinvlp_4
X_12325_ net646 net511 VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_11_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15113_ net956 net1026 _05043_ VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__and3_1
XFILLER_142_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16093_ _06956_ _06963_ _06964_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__nand3_1
XFILLER_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _09439_ _09646_ _03186_ _03187_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__o211ai_1
XFILLER_48_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19921_ _01135_ _01138_ _00994_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__nand3_4
X_15044_ net726 net723 net861 net668 VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__and4_1
X_11207_ net990 _02126_ net228 VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__a21oi_4
X_12187_ _03119_ _03117_ _03116_ VGND VGND VPWR VPWR _03122_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19852_ _01054_ _01056_ _01061_ _01062_ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__nand4_1
XFILLER_122_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11138_ _02006_ _02079_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__nand2_1
XFILLER_68_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18803_ _09694_ _09693_ VGND VGND VPWR VPWR _09696_ sky130_fd_sc_hd__nor2_1
X_16995_ _07703_ _07716_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__nand2_1
XFILLER_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19783_ net366 _00990_ _00987_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__and3_1
X_15946_ net261 _06821_ _06823_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__o21ai_1
X_11069_ _09428_ _09592_ net1062 _02007_ _02005_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__o221ai_2
X_18734_ _09614_ _09618_ _09598_ net335 VGND VGND VPWR VPWR _09620_ sky130_fd_sc_hd__o211a_1
XFILLER_48_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
X_15877_ net595 _06680_ net541 _06682_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__a31o_1
X_18665_ _09540_ _09541_ _09531_ VGND VGND VPWR VPWR _09545_ sky130_fd_sc_hd__and3_1
XFILLER_37_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17616_ net578 net479 VGND VGND VPWR VPWR _08480_ sky130_fd_sc_hd__nand2_1
X_14828_ _05726_ _05727_ _05714_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__a21oi_4
X_18596_ _09462_ _09464_ _09467_ VGND VGND VPWR VPWR _09469_ sky130_fd_sc_hd__a21oi_1
X_17547_ _08390_ _08405_ _08407_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__nand3_1
X_14759_ _05658_ _05659_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__nand2_1
X_17478_ _08187_ _08189_ _08191_ _08197_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__a31oi_1
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16429_ _07297_ _07298_ _07299_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__nand3_1
X_19217_ _10071_ _10110_ _10112_ VGND VGND VPWR VPWR _10114_ sky130_fd_sc_hd__nand3_4
XFILLER_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19148_ _09931_ _10034_ _10035_ _10037_ VGND VGND VPWR VPWR _10040_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_106_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19079_ _09968_ _09964_ _09967_ VGND VGND VPWR VPWR _09970_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_93_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20756_ clknet_leaf_52_clk _00396_ VGND VGND VPWR VPWR p_ll\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ _01595_ _01599_ net443 _01603_ _01605_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__a311o_1
X_20687_ clknet_3_0__leaf_clk _00327_ VGND VGND VPWR VPWR p_hl\[21\] sky130_fd_sc_hd__dfxtp_2
XFILLER_136_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10371_ _01354_ _01364_ _01268_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__nor3_1
XFILLER_123_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12110_ _03042_ _03044_ net706 net475 VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__and4_4
X_13090_ _09515_ _09657_ _03891_ _03963_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__o31a_1
XFILLER_2_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12041_ net658 net511 VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__nand2_4
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15800_ net602 net531 VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__nand2_1
X_16780_ _07644_ _07647_ _07640_ VGND VGND VPWR VPWR _07651_ sky130_fd_sc_hd__a21o_1
X_13992_ net788 net783 net650 net643 VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__nand4_2
X_15731_ net1070 _06605_ _06599_ _06604_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__o211ai_2
X_12943_ _03711_ _03783_ _03782_ VGND VGND VPWR VPWR _03871_ sky130_fd_sc_hd__a21boi_1
X_18450_ _09304_ _09306_ _09191_ VGND VGND VPWR VPWR _09311_ sky130_fd_sc_hd__a21o_1
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15662_ _06536_ _06537_ _06535_ VGND VGND VPWR VPWR _06543_ sky130_fd_sc_hd__a21oi_2
X_17401_ _08036_ _08038_ _08264_ _08265_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__nand4_2
X_12874_ _09460_ _09679_ _03799_ _03800_ VGND VGND VPWR VPWR _03802_ sky130_fd_sc_hd__o211ai_2
XFILLER_121_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11825_ _02648_ _02657_ _02659_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__o21ai_1
X_15593_ net612 net540 VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__nand2_1
X_18381_ net782 net584 VGND VGND VPWR VPWR _09235_ sky130_fd_sc_hd__nand2_1
XFILLER_61_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14613_ _05510_ _05512_ _05509_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11756_ _02679_ _02683_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__nand2_1
X_17332_ _08115_ _08119_ _08192_ _08194_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_16_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ net767 net1135 VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__nand2_4
X_17263_ _08124_ _08125_ net235 VGND VGND VPWR VPWR _08131_ sky130_fd_sc_hd__a21oi_1
X_10707_ _01739_ _01737_ _01736_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__a21o_1
XFILLER_41_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14475_ net193 _05375_ _05376_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__nand3_4
X_16214_ _07014_ _06974_ _07015_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__a21o_4
X_11687_ net325 _02624_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__nand2_1
X_13426_ net766 net689 VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__nand2_1
X_19002_ _09891_ _09884_ _09881_ _09892_ VGND VGND VPWR VPWR _09893_ sky130_fd_sc_hd__o211a_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10638_ _01676_ _01678_ _01681_ _01682_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__o2bb2ai_2
X_17194_ _08051_ _08057_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__nand2_1
X_16145_ _06974_ _07014_ _07016_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__nand3_2
X_13357_ _04241_ _04232_ _04230_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__a21o_1
X_10569_ net794 net1287 VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__and2_1
X_16076_ _06926_ _06932_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__nand2_1
X_12308_ _03238_ _03239_ _03240_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__a21o_1
XFILLER_127_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13288_ _04200_ _04201_ _04189_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__a21o_1
X_12239_ _02973_ _02981_ _02982_ _02990_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__a31oi_2
XFILLER_5_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15027_ net730 net663 VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__nand2_1
X_19904_ _01113_ _01122_ _01118_ _01123_ VGND VGND VPWR VPWR _01124_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_75_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19835_ _01040_ _01048_ _01046_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__o21ai_2
X_16978_ _07842_ _07843_ _07777_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__a21o_1
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19766_ _00713_ _00972_ _00971_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__a21oi_4
X_15929_ _06799_ _06800_ _06804_ VGND VGND VPWR VPWR _06807_ sky130_fd_sc_hd__nand3_2
Xinput4 a[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_18717_ _09533_ _09536_ _09539_ VGND VGND VPWR VPWR _09601_ sky130_fd_sc_hd__o21a_1
X_19697_ net591 net588 net729 net725 VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__and4_1
X_18648_ _09446_ _09523_ VGND VGND VPWR VPWR _09527_ sky130_fd_sc_hd__nand2_1
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18579_ net610 net749 VGND VGND VPWR VPWR _09451_ sky130_fd_sc_hd__and2_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20610_ clknet_leaf_35_clk _00250_ VGND VGND VPWR VPWR p_ll_pipe\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20541_ clknet_leaf_42_clk _00181_ VGND VGND VPWR VPWR mid_sum\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20472_ clknet_leaf_37_clk _00112_ VGND VGND VPWR VPWR term_mid\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_87_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _02473_ _02474_ _02546_ _02547_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__nand4_2
X_12590_ _03515_ _03519_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__nand2_1
XFILLER_70_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20808_ clknet_leaf_0_clk _00448_ VGND VGND VPWR VPWR b_h\[14\] sky130_fd_sc_hd__dfxtp_2
XFILLER_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11541_ _02366_ _02368_ _02355_ _02379_ _02381_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__a32oi_4
XTAP_TAPCELL_ROW_13_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ clknet_leaf_36_clk _00379_ VGND VGND VPWR VPWR p_ll\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire424 _05832_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_1
X_11472_ _02407_ _02409_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__nand2_1
Xwire435 _04323_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_1
XFILLER_7_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14260_ _05161_ _05163_ _09155_ _09515_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__o2bb2ai_1
Xwire446 _09799_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_2
X_10423_ _01574_ _01582_ _01585_ _01580_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__o211a_1
XFILLER_137_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13211_ _04129_ _04131_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__nor2_1
X_14191_ _04953_ _04957_ _05093_ _05094_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__a22oi_2
X_13142_ _04024_ _04027_ _04063_ _04064_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__nand4_1
X_10354_ term_low\[30\] term_mid\[30\] VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__xnor2_1
X_17950_ _08790_ _08801_ _08805_ net1104 VGND VGND VPWR VPWR _08807_ sky130_fd_sc_hd__o22ai_1
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13073_ _03998_ _03997_ net65 VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a21oi_1
X_10285_ _00504_ _00515_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__nor2_1
XFILLER_3_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12024_ _02590_ _02694_ _02955_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__o21ai_1
X_16901_ _07766_ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__nand2_1
X_17881_ _08737_ _08740_ _08739_ VGND VGND VPWR VPWR _08741_ sky130_fd_sc_hd__o21ai_1
X_16832_ _07556_ _07590_ _07699_ _07700_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__o211ai_4
Xclone303 net623 VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__clkbuf_16
Xclone314 net599 VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19620_ _00809_ _00813_ _00814_ _00782_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__o211ai_4
XFILLER_120_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19551_ b_l\[6\] net755 net562 net556 VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__and4_1
X_16763_ _06999_ _07632_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__or2_4
X_18502_ net459 _07100_ _09234_ VGND VGND VPWR VPWR _09367_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13975_ _09471_ _09482_ net805 _04874_ _04879_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__o311a_1
X_16694_ _07564_ _07565_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__nand2_1
X_15714_ _06588_ _06589_ _06587_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__a21oi_2
X_12926_ _03846_ _03808_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__nand2_1
XFILLER_19_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19482_ _00661_ _00662_ _00665_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__a21oi_1
X_15645_ _06525_ _06517_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__nand2_1
X_12857_ _03781_ _03784_ _03785_ _03709_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__o211ai_4
X_18433_ _09265_ _09266_ _09289_ VGND VGND VPWR VPWR _09292_ sky130_fd_sc_hd__nand3_1
XFILLER_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11808_ _02740_ _02736_ _02732_ _02741_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__o211ai_2
X_18364_ net626 net737 VGND VGND VPWR VPWR _09216_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_32_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15576_ _06454_ _06427_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__nand2_1
X_17315_ net585 net485 net479 net593 VGND VGND VPWR VPWR _08182_ sky130_fd_sc_hd__a22o_1
X_12788_ net680 _03629_ net475 _03627_ VGND VGND VPWR VPWR _03717_ sky130_fd_sc_hd__a31o_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11739_ _02673_ _02572_ _02674_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__nand3_2
X_18295_ _09136_ _09138_ _09134_ VGND VGND VPWR VPWR _09141_ sky130_fd_sc_hd__a21oi_1
X_14527_ _05417_ _05423_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__nand2_2
X_17246_ _08110_ _08107_ _08103_ _08111_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__o211ai_2
X_14458_ _05360_ _05137_ _05359_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__and3_1
Xmax_cap702 net706 VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__buf_6
X_17177_ _08043_ _08044_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13409_ _04303_ _04268_ _04301_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a21oi_2
X_14389_ _05277_ _05279_ _05288_ _05289_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__nand4_2
X_16128_ _06996_ _06997_ _06995_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__o21ai_1
Xmax_cap713 a_h\[0\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__buf_8
Xmax_cap746 net748 VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__buf_12
Xmax_cap735 net915 VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__buf_8
Xmax_cap779 net780 VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__buf_8
Xmax_cap768 net770 VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__buf_12
Xmax_cap757 net758 VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__buf_12
X_16059_ _06846_ _06930_ _06931_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__nand3b_4
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19818_ _01031_ _01012_ VGND VGND VPWR VPWR _01032_ sky130_fd_sc_hd__nand2_1
XFILLER_29_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19749_ _00867_ _00953_ _00955_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__nand3_1
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_31 _00050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _01860_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20524_ clknet_leaf_43_clk _00164_ VGND VGND VPWR VPWR term_low\[19\] sky130_fd_sc_hd__dfxtp_1
X_20455_ clknet_leaf_16_clk _00095_ VGND VGND VPWR VPWR term_high\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20386_ clknet_leaf_41_clk _00026_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfxtp_1
XFILLER_121_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10972_ net691 net538 VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__nand2_1
X_13760_ _04665_ net432 _04556_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__o21ai_2
XFILLER_71_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12711_ net648 b_h\[9\] net829 net1015 VGND VGND VPWR VPWR _03641_ sky130_fd_sc_hd__a22oi_1
X_13691_ _09155_ _09471_ _02362_ _04134_ _04596_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__o221a_1
X_12642_ _03534_ _03571_ _03572_ VGND VGND VPWR VPWR _03573_ sky130_fd_sc_hd__nand3_2
X_15430_ _06320_ _06321_ net716 net650 VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__nand4_1
XFILLER_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12573_ _03415_ net246 _03456_ _03455_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__a31o_1
X_15361_ _06253_ _06254_ _06220_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__a21oi_2
XFILLER_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11524_ _02450_ _02457_ _02458_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__nand3_1
X_17100_ net612 net476 _07968_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__a21oi_1
X_18080_ _08915_ _08925_ _08926_ VGND VGND VPWR VPWR _08929_ sky130_fd_sc_hd__nand3_4
Xwire232 _09181_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
X_14312_ _05213_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nand2_1
Xwire210 _05083_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_1
X_15292_ _06185_ _06186_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__nand2_2
X_11455_ net1078 net510 VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__nand2_1
X_17031_ _07642_ net530 net550 VGND VGND VPWR VPWR _07900_ sky130_fd_sc_hd__nand3_1
XFILLER_8_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14243_ net761 net662 VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__nand2_1
X_10406_ _01575_ _01576_ _01577_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__a21boi_2
XFILLER_137_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire298 _00451_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_4
X_11386_ _02240_ _02319_ _02320_ _02223_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a31o_1
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14174_ _05075_ net316 VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__nand2_1
X_13125_ _04047_ _04048_ VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__or2_1
X_18982_ net618 net729 net725 net621 VGND VGND VPWR VPWR _09873_ sky130_fd_sc_hd__a22o_4
X_10337_ term_low\[28\] term_mid\[28\] VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nor2_1
X_17933_ _08788_ _08789_ VGND VGND VPWR VPWR _08791_ sky130_fd_sc_hd__nand2b_1
X_10268_ term_low\[17\] term_mid\[17\] VGND VGND VPWR VPWR _10072_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _03923_ _03978_ _03980_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__nand3_1
X_12007_ net247 _02942_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__nor2_1
XFILLER_94_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17864_ _08722_ _08723_ VGND VGND VPWR VPWR _08724_ sky130_fd_sc_hd__xnor2_1
X_19603_ net579 net836 net574 net918 VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__nand4_4
X_10199_ net722 VGND VGND VPWR VPWR _09351_ sky130_fd_sc_hd__inv_6
X_16815_ _07678_ _07683_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__nand2_1
X_17795_ _08655_ _08656_ _08646_ VGND VGND VPWR VPWR _08657_ sky130_fd_sc_hd__a21o_1
Xclone166 a_h\[1\] VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__clkbuf_16
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16746_ _07614_ _07615_ _07599_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__a21o_1
X_19534_ _00724_ _00725_ _00722_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__a21o_1
X_13958_ _04856_ _04857_ _04860_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__nand3_1
X_12909_ _03821_ _03833_ _03834_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__nand3_2
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19465_ net755 net567 net562 net879 VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__a22o_1
X_16677_ _07509_ _07546_ _07547_ VGND VGND VPWR VPWR _07549_ sky130_fd_sc_hd__nand3_2
X_18416_ net610 net759 net754 net802 VGND VGND VPWR VPWR _09273_ sky130_fd_sc_hd__a22oi_1
X_13889_ _04788_ _04791_ net714 net728 VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__nand4_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15628_ _06506_ net512 net632 VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__nand3_2
X_19396_ _00537_ _00543_ _00555_ _00541_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__o22ai_2
X_15559_ net625 net628 net532 net528 VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__nand4_2
X_18347_ _09182_ _09185_ net276 _09192_ VGND VGND VPWR VPWR _09198_ sky130_fd_sc_hd__o2bb2ai_1
X_18278_ _09114_ _09122_ _09123_ VGND VGND VPWR VPWR _09124_ sky130_fd_sc_hd__nand3_4
XFILLER_30_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17229_ net600 net593 net485 net479 VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__nand4_2
Xinput40 b[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap521 net523 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_12
Xmax_cap510 net511 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_12
Xinput51 b[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput62 b[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
Xmax_cap543 net544 VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__buf_12
Xmax_cap532 net533 VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__buf_8
Xmax_cap554 net555 VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_12
X_20240_ _01480_ _01481_ net250 VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__nand3_1
Xmax_cap587 net590 VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_114_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap565 net566 VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__buf_12
Xmax_cap576 net577 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__buf_8
X_20171_ net724 net551 VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__nand2_2
Xmax_cap598 net599 VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__buf_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20507_ clknet_leaf_35_clk _00147_ VGND VGND VPWR VPWR term_low\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_5_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20438_ clknet_leaf_13_clk _00078_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfxtp_1
X_11240_ _02178_ _02163_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__nand2_2
X_11171_ _02103_ _02112_ _02113_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__nand3b_1
XFILLER_107_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20369_ clknet_leaf_48_clk _00009_ VGND VGND VPWR VPWR b_l\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_106_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14930_ _05824_ _05825_ _05826_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_145_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14861_ net715 net1009 _05754_ _05755_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__a22o_4
X_16600_ a_l\[2\] net620 net484 net480 VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__and4_1
XFILLER_91_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17580_ _08429_ _08431_ _08443_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_3_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13812_ _04608_ _04703_ _04712_ _04713_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__o211ai_2
X_16531_ net307 _07389_ _07396_ _07397_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_90_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14792_ _05689_ _05678_ _05688_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__nand3_2
X_10955_ _01900_ _01901_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__nand2_1
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13743_ _04625_ net287 _04647_ _04648_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_43_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16462_ _07330_ _07332_ _07320_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__o21ai_1
X_13674_ _04485_ _04580_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__nand2_1
X_10886_ net794 net1253 VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__and2_1
X_19250_ _09991_ _09736_ _09994_ VGND VGND VPWR VPWR _10151_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16393_ _07261_ _07263_ net930 net502 VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__nand4_4
X_12625_ _03551_ _03552_ _03553_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__a21o_1
X_18201_ net800 net764 VGND VGND VPWR VPWR _09048_ sky130_fd_sc_hd__nand2_1
X_15413_ _06217_ _06303_ _06305_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_42_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19181_ _09917_ _09920_ _09918_ VGND VGND VPWR VPWR _10076_ sky130_fd_sc_hd__a21boi_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12556_ _03483_ _03486_ _03377_ VGND VGND VPWR VPWR _03488_ sky130_fd_sc_hd__o21ai_2
X_18132_ _08975_ _08976_ _08979_ VGND VGND VPWR VPWR _08980_ sky130_fd_sc_hd__nand3_4
X_15344_ _06237_ _06236_ _06235_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_42_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _02247_ _02431_ _02430_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__o21ai_1
XFILLER_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18063_ _08905_ _08906_ _08911_ VGND VGND VPWR VPWR _08912_ sky130_fd_sc_hd__a21oi_1
X_12487_ net633 net518 VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__and2_1
X_15275_ _06163_ _06166_ _09308_ _09515_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_137_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17014_ _07882_ _07883_ net796 VGND VGND VPWR VPWR _07884_ sky130_fd_sc_hd__a21oi_1
X_11438_ _02376_ _02377_ _09439_ _09602_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__o2bb2a_1
X_14226_ _05125_ _05128_ _05122_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__a21o_1
X_11369_ _02303_ _02273_ _02304_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__nand3_4
XFILLER_98_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14157_ _05055_ _05058_ _05052_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__a21o_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13108_ _04030_ _04032_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__nand2_2
X_18965_ _09716_ _09722_ _09854_ _09855_ VGND VGND VPWR VPWR _09857_ sky130_fd_sc_hd__a22oi_1
X_14088_ _04981_ _04992_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__nand2_2
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17916_ _08709_ _08743_ _08771_ _08714_ _08744_ VGND VGND VPWR VPWR _08775_ sky130_fd_sc_hd__a221o_1
X_13039_ net1049 net634 net826 net885 VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__and4_1
X_18896_ _09680_ _09683_ _09685_ VGND VGND VPWR VPWR _09788_ sky130_fd_sc_hd__o21ai_2
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17847_ _08706_ _08707_ _08662_ VGND VGND VPWR VPWR _08708_ sky130_fd_sc_hd__nand3_1
XFILLER_66_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17778_ _08494_ _08635_ _08636_ _08634_ VGND VGND VPWR VPWR _08640_ sky130_fd_sc_hd__o211ai_2
X_19517_ net1080 _00576_ _00705_ _00706_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__nand4_4
X_16729_ _07455_ _07458_ _07460_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__o21ai_1
X_19448_ _00628_ _00630_ _00589_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__nand3_2
X_19379_ _00542_ _00544_ _00554_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_116_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer217 net710 VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_20_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer206 _00682_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__buf_2
Xrebuffer228 a_h\[10\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap362 _02163_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
Xmax_cap340 _08313_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_4
X_20223_ _01458_ _01465_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__nand2_1
XFILLER_143_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap384 net387 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
Xmax_cap373 _08960_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
Xmax_cap395 _03909_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_2
X_20154_ net215 net251 _01389_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__nand3_2
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20085_ _01315_ _01316_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__a21o_1
XFILLER_85_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ p_hl\[17\] p_lh\[17\] _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__o21ai_1
X_10671_ _09537_ _09548_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o21ai_1
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12410_ _03295_ _03298_ _03337_ _03339_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__nand4_2
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13390_ _04299_ _04293_ _04270_ _04300_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__o211ai_2
XFILLER_139_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12341_ _03268_ _03269_ _03253_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__and3_1
XFILLER_5_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12272_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__nand3_1
X_15060_ _05955_ _05957_ _05919_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__a21o_1
X_11223_ net1061 net536 VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__nand2_1
X_14011_ _04913_ _04916_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__nand2_1
XFILLER_122_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ _02086_ _02090_ _02092_ _02073_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__o211ai_1
XFILLER_108_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11085_ _02015_ _02017_ _02026_ _02027_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__o2bb2ai_2
X_15962_ _06837_ _06838_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__nand2_1
XFILLER_95_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18750_ net301 _09508_ _09496_ VGND VGND VPWR VPWR _09638_ sky130_fd_sc_hd__a21boi_1
X_17701_ net555 net940 net500 net494 VGND VGND VPWR VPWR _08564_ sky130_fd_sc_hd__nand4_4
XFILLER_76_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18681_ _09529_ _09530_ _09557_ _09560_ VGND VGND VPWR VPWR _09563_ sky130_fd_sc_hd__o2bb2ai_4
X_14913_ _05806_ _05808_ _05809_ VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__a21o_1
X_15893_ net613 net515 VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__nand2_1
XFILLER_75_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17632_ _08490_ _08491_ _08494_ _08395_ VGND VGND VPWR VPWR _08496_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_75_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14844_ _05740_ _05742_ _05708_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__o21ai_4
X_11987_ _02910_ _02915_ _02917_ _02880_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__o211ai_2
X_17563_ _08420_ _08414_ _08382_ _08419_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_67_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14775_ net767 net761 net640 net636 VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__and4_1
X_10938_ net702 net1106 VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__nand2_1
X_16514_ _07375_ _07383_ _07385_ _07384_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__o211ai_2
X_17494_ _08357_ _08341_ _08284_ _08358_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__o211ai_2
X_19302_ net984 _00469_ _00470_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__a21oi_1
X_13726_ net751 net694 net689 net757 VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__a22o_1
XFILLER_140_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16445_ _09166_ _09668_ _02589_ _06441_ _07314_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__o221a_1
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19233_ _10128_ _10130_ VGND VGND VPWR VPWR _10132_ sky130_fd_sc_hd__nor2_2
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10869_ net793 net1318 VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__and2_1
XFILLER_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13657_ _04553_ _04551_ _04561_ net264 VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__o2bb2ai_4
X_16376_ _07243_ _07245_ net587 net515 VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__and4_1
X_12608_ net659 net980 net995 net495 VGND VGND VPWR VPWR _03539_ sky130_fd_sc_hd__nand4_4
X_13588_ _04401_ _04404_ _04405_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19164_ _10039_ _10040_ _10048_ _10051_ VGND VGND VPWR VPWR _10057_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_144_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12539_ _03331_ _03467_ _03468_ _03466_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__a31oi_1
X_18115_ _08913_ _08929_ _08927_ _08922_ VGND VGND VPWR VPWR _08963_ sky130_fd_sc_hd__o2bb2ai_4
X_19095_ _09979_ _09981_ net630 net717 VGND VGND VPWR VPWR _09986_ sky130_fd_sc_hd__nand4_1
X_15327_ net726 net643 VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__nand2_2
X_18046_ net630 net759 VGND VGND VPWR VPWR _08895_ sky130_fd_sc_hd__nand2_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15258_ _09362_ _09482_ _06149_ _06151_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__o22a_1
XFILLER_144_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14209_ _09177_ _09384_ _05109_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__o21a_1
X_15189_ _06010_ _06012_ _06037_ _06041_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__o211ai_2
XFILLER_141_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19997_ _01220_ _01221_ _01110_ _01218_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__o2bb2ai_1
X_18948_ _09794_ _09835_ _09837_ VGND VGND VPWR VPWR _09840_ sky130_fd_sc_hd__and3_1
XFILLER_104_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_66_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18879_ _09769_ _09770_ VGND VGND VPWR VPWR _09771_ sky130_fd_sc_hd__nand2_4
XFILLER_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20772_ clknet_leaf_0_clk _00412_ VGND VGND VPWR VPWR a_h\[10\] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold440 p_hh_pipe\[17\] VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap170 _08799_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
Xhold462 mid_sum\[2\] VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 p_ll_pipe\[28\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold495 p_hh_pipe\[7\] VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 p_hh_pipe\[24\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 p_hh_pipe\[25\] VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap192 _06359_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
Xmax_cap181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
X_20206_ _01396_ _01398_ _01445_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20137_ net568 net721 _01371_ _01372_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__a22o_1
XFILLER_100_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20068_ net742 net735 net551 net549 _01293_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_142_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _02843_ _02845_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__nand2_1
X_12890_ _03814_ _03816_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__nor2_1
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11841_ _09406_ _09646_ _02773_ _02775_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_107_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ net679 net1048 net511 net508 VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__nand4_1
X_14560_ _05455_ _05457_ _05437_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__o21ai_2
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10723_ _01747_ _01751_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__and2_1
X_13511_ _09155_ _09449_ _04349_ _04416_ _04415_ VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_49_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14491_ _05393_ _05392_ _05267_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__nand3_4
X_16230_ _09592_ _07101_ _07094_ _07099_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__o211a_1
X_10654_ p_hl\[4\] p_lh\[4\] _01687_ _01690_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__o22ai_1
XTAP_TAPCELL_ROW_62_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13442_ net777 net935 _04351_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a22oi_4
X_16161_ _07035_ _07036_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__nor2_2
X_10585_ net793 net1225 VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__and2_1
X_13373_ net785 net934 net675 net787 VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__a22oi_4
Xclkload29 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__inv_4
X_12324_ net1019 b_h\[8\] VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__nand2_1
XFILLER_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload18 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_8
XFILLER_5_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15112_ net722 net661 VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__nand2_1
X_16092_ _06955_ _06965_ _06966_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__nand3_1
XFILLER_127_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12255_ _03186_ _03187_ _03188_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__a21o_1
X_19920_ _00993_ _00985_ _01141_ _01140_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__o211ai_4
X_15043_ net726 net668 VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__nand2_1
X_11206_ _02139_ _02147_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__nor2_1
X_12186_ _03120_ _02959_ _02818_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__nand3_2
X_19851_ _00954_ _00867_ _00953_ _01066_ _01067_ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__o2111ai_4
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11137_ net671 net965 net538 net1061 VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__a22oi_4
X_18802_ _09693_ _09694_ VGND VGND VPWR VPWR _09695_ sky130_fd_sc_hd__and2_1
X_19782_ _00990_ _00987_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__nand2_1
X_16994_ _07850_ _07852_ _07858_ _07859_ VGND VGND VPWR VPWR _07864_ sky130_fd_sc_hd__nand4_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18733_ _09617_ net447 _09601_ _09615_ VGND VGND VPWR VPWR _09619_ sky130_fd_sc_hd__o211ai_2
X_15945_ _06749_ _06819_ _06820_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__nand3_4
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11068_ net1062 _02007_ net967 net1106 _02005_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__o2111ai_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15876_ _06680_ _06753_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__nand2_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18664_ _09532_ _09542_ _09543_ VGND VGND VPWR VPWR _09544_ sky130_fd_sc_hd__nand3_2
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17615_ _08210_ net503 net550 VGND VGND VPWR VPWR _08479_ sky130_fd_sc_hd__and3_1
X_18595_ _09462_ _09464_ _09467_ VGND VGND VPWR VPWR _09468_ sky130_fd_sc_hd__and3_1
X_14827_ _05722_ _05723_ _05725_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__nand3_4
X_17546_ _08405_ _08407_ _08390_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__a21o_1
X_14758_ _05654_ _05653_ _05537_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__nand3_2
X_17477_ _08182_ net476 net600 _08180_ VGND VGND VPWR VPWR _08343_ sky130_fd_sc_hd__a31o_1
X_13709_ net456 _04613_ _04616_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__o21ai_2
X_14689_ _05561_ net312 _05587_ _05588_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__nand4_2
X_16428_ _07297_ _07298_ _07299_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__and3_1
X_19216_ _10070_ _10071_ _10109_ _10111_ VGND VGND VPWR VPWR _10113_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_4_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16359_ _07230_ _07231_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__nand2_2
X_19147_ _09931_ _10034_ _10036_ _10038_ VGND VGND VPWR VPWR _10039_ sky130_fd_sc_hd__nand4_4
XFILLER_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19078_ _09960_ _09924_ _09835_ _09963_ VGND VGND VPWR VPWR _09969_ sky130_fd_sc_hd__a22oi_2
XFILLER_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18029_ _08876_ _08867_ _08875_ VGND VGND VPWR VPWR _08879_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_93_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20755_ clknet_leaf_49_clk _00395_ VGND VGND VPWR VPWR p_ll\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20686_ clknet_leaf_57_clk _00326_ VGND VGND VPWR VPWR p_hl\[20\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_102_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10370_ term_low\[31\] term_mid\[31\] _01428_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__a21o_1
XFILLER_105_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ net1048 net501 VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13991_ net788 net783 net650 VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__nand3_1
X_15730_ net966 net541 _06604_ _06607_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__a22o_1
X_12942_ _03862_ _03866_ _03868_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__and3_1
XFILLER_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15661_ _06539_ _06540_ _06534_ VGND VGND VPWR VPWR _06542_ sky130_fd_sc_hd__a21o_1
XFILLER_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17400_ _08264_ _08265_ _08266_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__a21bo_1
X_12873_ net674 net473 VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__nand2_1
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14612_ _09384_ _09395_ _05510_ _05512_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__o211ai_1
XFILLER_27_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11824_ net248 _02760_ _02759_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__o21ai_1
X_15592_ _06439_ _06437_ _06442_ VGND VGND VPWR VPWR _06474_ sky130_fd_sc_hd__a21bo_1
X_18380_ net780 net585 VGND VGND VPWR VPWR _09234_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _02571_ _02691_ _02692_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__o21a_1
X_17331_ _08115_ _08119_ _08192_ _08194_ VGND VGND VPWR VPWR _08198_ sky130_fd_sc_hd__o22a_1
XFILLER_14_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _05442_ _05443_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__nand2_1
X_17262_ _07963_ _08088_ _08123_ _08124_ VGND VGND VPWR VPWR _08130_ sky130_fd_sc_hd__a22o_1
X_10706_ _01737_ _01739_ _01741_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__o21a_1
XFILLER_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14474_ _05268_ _05374_ _05373_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nand3_4
X_16213_ _07086_ _07087_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__nand2_2
X_11686_ _02619_ _02618_ _02621_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__nand3_4
X_13425_ net763 net701 VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nand2_1
X_19001_ _09885_ _09886_ _09199_ _09308_ VGND VGND VPWR VPWR _09892_ sky130_fd_sc_hd__o2bb2ai_1
X_10637_ _01681_ _01682_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__nor2_1
X_17193_ _08054_ _08057_ _08051_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__a21o_1
X_16144_ _07014_ _07016_ _06974_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13356_ _04266_ _04267_ VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__and2_4
X_10568_ net794 net1298 VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__and2_1
X_10499_ _01653_ term_high\[52\] net1331 VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__a21oi_1
X_16075_ _06927_ net238 _06925_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__a21oi_2
X_12307_ _03238_ _03239_ _03240_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__a21oi_1
X_13287_ _04163_ _04190_ _04198_ _04199_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__o211ai_2
XFILLER_5_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12238_ _03169_ _03171_ VGND VGND VPWR VPWR _03172_ sky130_fd_sc_hd__nand2_1
X_15026_ _05826_ _05823_ _05825_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__o21ai_1
X_19903_ _01112_ _01114_ _01109_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__a21o_1
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12169_ _02967_ _03099_ _03100_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__nand3_1
XFILLER_110_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19834_ _01001_ _01041_ _01043_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__nand3_1
X_16977_ _07773_ _07774_ _07842_ _07843_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__a22oi_2
XFILLER_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19765_ _10004_ _00974_ _10002_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__nand3_4
X_15928_ _06801_ _06802_ _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__nand3_2
XFILLER_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput5 a[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18716_ _09533_ _09536_ _09539_ VGND VGND VPWR VPWR _09600_ sky130_fd_sc_hd__o21ai_1
X_19696_ net588 net729 VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__nand2_1
X_18647_ _09514_ _09517_ _09473_ _09512_ VGND VGND VPWR VPWR _09525_ sky130_fd_sc_hd__o211ai_4
X_15859_ _06734_ _06735_ _06737_ _06650_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__o2bb2ai_4
X_18578_ _09357_ _09447_ VGND VGND VPWR VPWR _09450_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_35_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17529_ a_l\[11\] net488 VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__nand2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20540_ clknet_leaf_42_clk net365 VGND VGND VPWR VPWR mid_sum\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20471_ clknet_leaf_12_clk _00111_ VGND VGND VPWR VPWR term_high\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_114_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_67_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20807_ clknet_leaf_4_clk _00447_ VGND VGND VPWR VPWR b_h\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11540_ _02389_ _02477_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__nand2_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire403 _02024_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__buf_1
X_20738_ clknet_leaf_35_clk _00378_ VGND VGND VPWR VPWR p_ll\[8\] sky130_fd_sc_hd__dfxtp_1
Xwire414 _08472_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_567 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11471_ _02407_ _02408_ _02409_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__a21o_1
Xwire436 _03546_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_1
X_20669_ clknet_leaf_5_clk _00309_ VGND VGND VPWR VPWR p_hl\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10422_ _01565_ _01575_ _01580_ _01585_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__and4_1
Xwire469 _01717_ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_1
X_13210_ net793 _04128_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__nand2_1
X_14190_ _04953_ _04957_ _05093_ _05094_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__nand4_1
XFILLER_124_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13141_ _04024_ _04027_ _04063_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a22oi_1
X_10353_ net1368 term_mid\[30\] VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_76_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13072_ _03956_ _03948_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__nand2_1
X_12023_ _02953_ _02957_ _02810_ _02958_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__o211ai_4
X_16900_ _07767_ _07769_ _07736_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__nand3_4
X_10284_ _10148_ _10169_ _00493_ net797 VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__a31o_1
X_17880_ _08699_ _08735_ _08738_ VGND VGND VPWR VPWR _08740_ sky130_fd_sc_hd__a21o_1
X_16831_ _07696_ _07697_ _07628_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__a21o_1
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16762_ net571 net566 net523 net516 VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__and4_1
XFILLER_76_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19550_ net880 net556 VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__nand2_1
XFILLER_19_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15713_ net624 net515 _06592_ _06591_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__a22oi_4
X_18501_ net459 _07100_ _09234_ VGND VGND VPWR VPWR _09366_ sky130_fd_sc_hd__o21a_1
X_13974_ _04876_ _04878_ net762 net670 VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__o211a_1
X_16693_ _07559_ _07451_ _07558_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__nand3_4
XPHY_EDGE_ROW_85_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12925_ _03809_ _03844_ _03845_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__nand3_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19481_ _00661_ _00662_ _00664_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__nand3_2
X_15644_ _06440_ _06521_ _06524_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__o21ai_1
X_12856_ _03782_ _03783_ _03711_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__a21o_1
X_18432_ _09265_ _09289_ VGND VGND VPWR VPWR _09291_ sky130_fd_sc_hd__nand2_1
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15575_ _06425_ _06454_ _06455_ _06410_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__and4_1
X_11807_ _02740_ _02736_ _02732_ _02741_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__o211a_1
X_18363_ _09183_ _09176_ _09182_ _09195_ VGND VGND VPWR VPWR _09215_ sky130_fd_sc_hd__a22oi_2
XFILLER_33_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17314_ net585 net485 net479 net593 VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__a22oi_2
X_12787_ _09449_ _09679_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__nor2_1
X_14526_ _05427_ _05416_ _05426_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_32_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _02604_ _02670_ _02672_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__nand3b_1
X_18294_ _09199_ _09220_ net922 _06681_ _09138_ VGND VGND VPWR VPWR _09140_ sky130_fd_sc_hd__o221a_1
XFILLER_41_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11669_ net652 net535 VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__and2_1
X_17245_ _02338_ _07100_ net585 net488 _08108_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__o2111ai_4
X_14457_ _05337_ _05339_ net349 _05354_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__a22o_1
X_17176_ net550 net1023 net516 net554 VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _04268_ _04303_ _04301_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__a21o_1
Xmax_cap703 net705 VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__clkbuf_8
X_14388_ _05277_ _05279_ _05289_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__nand3_1
X_16127_ _06998_ _07001_ net966 net515 VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_94_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13339_ _04204_ _04208_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__nand2_1
Xmax_cap714 a_h\[0\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__buf_8
XFILLER_6_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap736 net915 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__buf_8
Xmax_cap725 net1095 VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__clkbuf_8
Xmax_cap769 net770 VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__buf_8
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap747 net748 VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__buf_6
Xmax_cap758 net760 VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__buf_8
XFILLER_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16058_ _06846_ _06929_ _06931_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_90_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15009_ net756 net750 net640 net635 VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__nand4_4
XFILLER_110_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19817_ _01028_ _01030_ VGND VGND VPWR VPWR _01031_ sky130_fd_sc_hd__nand2_1
XFILLER_84_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19748_ _00953_ _00955_ _00867_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19679_ _00878_ _00880_ _00734_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__a21oi_2
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 _00434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _00350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20523_ clknet_leaf_42_clk _00163_ VGND VGND VPWR VPWR term_low\[18\] sky130_fd_sc_hd__dfxtp_1
X_20454_ clknet_leaf_16_clk _00094_ VGND VGND VPWR VPWR term_high\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20385_ clknet_leaf_31_clk _00025_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10971_ net697 net534 VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__nand2_1
XFILLER_90_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12710_ net1015 net976 net859 net830 VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__nand4_1
X_13690_ _02362_ _04134_ _04596_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__o21ai_1
XFILLER_43_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ _03395_ _03407_ _03563_ _03565_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__a22o_1
XFILLER_70_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12572_ _03415_ net246 _03456_ _03455_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__a31oi_4
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15360_ _06249_ _06251_ _06252_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__nand3b_4
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11523_ _02450_ _02457_ _02458_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__and3_1
XFILLER_8_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14311_ _05212_ _05202_ _05211_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__nand3_2
X_15291_ net284 _06182_ _06184_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__nand3_4
Xwire255 _07406_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__buf_1
X_11454_ net698 net501 VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__nand2_1
X_17030_ net554 net1038 _07811_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14242_ _04990_ _04993_ _04997_ net392 VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__a2bb2oi_2
Xwire244 _05036_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_1
X_10405_ _01575_ _01576_ net793 VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_59_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11385_ _02322_ _02323_ _02223_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__a21bo_1
XFILLER_124_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14173_ _05073_ _05074_ net316 VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__and3_1
X_13124_ _03966_ _04009_ _04046_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__and3_1
X_18981_ _09787_ _09788_ _09785_ VGND VGND VPWR VPWR _09872_ sky130_fd_sc_hd__a21oi_2
X_10336_ _01042_ _01053_ _01064_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__o21a_1
XFILLER_105_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17932_ _08789_ VGND VGND VPWR VPWR _08790_ sky130_fd_sc_hd__inv_2
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10267_ term_low\[17\] term_mid\[17\] VGND VGND VPWR VPWR _10061_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _03922_ _03979_ _03978_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__o21bai_2
X_12006_ _02789_ _02938_ _02939_ net474 net712 VGND VGND VPWR VPWR _02942_ sky130_fd_sc_hd__a32o_1
XFILLER_79_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17863_ _08494_ _08635_ _08685_ VGND VGND VPWR VPWR _08723_ sky130_fd_sc_hd__o21ai_2
XFILLER_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10198_ net560 VGND VGND VPWR VPWR _09340_ sky130_fd_sc_hd__clkinv_8
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19602_ _00797_ _00798_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__nand2_1
X_16814_ _07678_ _07681_ _07682_ _07496_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__o2bb2ai_2
X_17794_ a_l\[10\] net472 _08652_ _08653_ VGND VGND VPWR VPWR _08656_ sky130_fd_sc_hd__a22o_1
XFILLER_16_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone178 net499 VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__clkbuf_16
X_16745_ _07599_ _07614_ _07615_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__nand3_1
Xclone167 b_h\[6\] VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__clkbuf_16
X_19533_ _00615_ _00620_ _00630_ _00632_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__o211ai_4
X_13957_ _04858_ _04859_ _04861_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__nand3_1
X_16676_ _07540_ _07541_ _07510_ _07508_ net846 VGND VGND VPWR VPWR _07548_ sky130_fd_sc_hd__a32oi_4
XFILLER_62_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12908_ _03831_ _03832_ _03820_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__nand3_2
X_19464_ net755 net567 net562 b_l\[6\] VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__a22oi_2
X_15627_ _06506_ net512 net632 VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__and3_1
X_18415_ net610 net759 VGND VGND VPWR VPWR _09272_ sky130_fd_sc_hd__nand2_1
X_13888_ net714 net728 _04788_ _04791_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a22o_1
XFILLER_34_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12839_ _03654_ _03764_ net267 VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__o21ai_1
X_19395_ _10159_ _00560_ _00559_ _00563_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__a31o_1
XFILLER_15_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18346_ net276 _09192_ _09182_ _09185_ VGND VGND VPWR VPWR _09197_ sky130_fd_sc_hd__o211ai_1
X_15558_ net622 net888 VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__nand2_8
X_18277_ _09119_ net749 net626 _09118_ VGND VGND VPWR VPWR _09123_ sky130_fd_sc_hd__nand4_4
X_14509_ net193 _05375_ _05376_ _05377_ _05391_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__a32oi_4
X_15489_ _06376_ _06368_ _06375_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__or3_1
XFILLER_147_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput30 a[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_17228_ net600 net593 net485 net479 VGND VGND VPWR VPWR _08096_ sky130_fd_sc_hd__and4_1
Xmax_cap511 net514 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_12
Xmax_cap500 b_h\[9\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_12
Xinput52 b[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput41 b[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput63 b[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
X_17159_ _07584_ _07586_ _08024_ _08027_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__a31o_1
Xmax_cap544 net545 VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__buf_12
Xmax_cap522 net523 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_8
Xmax_cap533 net534 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_12
XFILLER_143_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_114_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap555 a_l\[14\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__buf_8
Xmax_cap566 a_l\[12\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__buf_12
Xmax_cap577 net578 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__buf_8
X_20170_ _01218_ net549 net731 VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__and3_1
Xmax_cap588 net589 VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__buf_12
XFILLER_143_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap599 net601 VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__buf_12
XFILLER_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20506_ clknet_leaf_35_clk _00146_ VGND VGND VPWR VPWR term_low\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20437_ clknet_leaf_13_clk _00077_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfxtp_1
X_11170_ _02106_ _02108_ _02109_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__a21o_1
X_20368_ clknet_leaf_48_clk _00008_ VGND VGND VPWR VPWR b_l\[8\] sky130_fd_sc_hd__dfxtp_4
XFILLER_134_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20299_ net551 b_l\[14\] net548 net716 _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__a41o_1
XFILLER_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14860_ _05754_ _05755_ net715 net1010 VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_3_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14791_ _05689_ _05678_ _05688_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__and3_1
X_13811_ _04714_ _04717_ _04705_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a21oi_2
X_16530_ _07391_ _07395_ _07398_ _07389_ net307 VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__o2111ai_2
XFILLER_113_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13742_ _04619_ _04624_ net287 _04649_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__o211ai_2
XFILLER_29_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10954_ _01875_ _01879_ _01898_ _01899_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a22o_1
XFILLER_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16461_ _07318_ _07319_ _07331_ _07333_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__o211ai_1
X_18200_ _08994_ _08980_ _08972_ _08981_ VGND VGND VPWR VPWR _09047_ sky130_fd_sc_hd__o2bb2ai_2
X_10885_ net794 net1294 VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__and2_1
XFILLER_71_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13673_ _04580_ _04581_ _04485_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__a21o_1
X_16392_ _09210_ _09613_ _07264_ _07265_ VGND VGND VPWR VPWR _07266_ sky130_fd_sc_hd__o211ai_4
X_12624_ _09439_ _09668_ _03551_ _03552_ VGND VGND VPWR VPWR _03555_ sky130_fd_sc_hd__o211ai_2
X_15412_ _06257_ net150 _06210_ _06258_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__a22oi_4
X_19180_ net1101 _09921_ VGND VGND VPWR VPWR _10075_ sky130_fd_sc_hd__nand2_1
X_12555_ net176 _03485_ _03484_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__o21ai_1
X_18131_ _08920_ _08977_ VGND VGND VPWR VPWR _08979_ sky130_fd_sc_hd__nand2_1
X_15343_ _06167_ _06171_ _06158_ _06174_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_42_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _02242_ _02243_ _02245_ _02430_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o31a_1
X_18062_ _08909_ net764 net627 VGND VGND VPWR VPWR _08911_ sky130_fd_sc_hd__nand3_1
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17013_ _07587_ _07728_ _07729_ _07726_ VGND VGND VPWR VPWR _07883_ sky130_fd_sc_hd__o2bb2a_1
X_12486_ _03415_ _03417_ VGND VGND VPWR VPWR _03418_ sky130_fd_sc_hd__nand2_1
X_15274_ _06163_ _06166_ _06160_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__a21oi_1
X_11437_ net678 net672 net525 net520 VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__nand4_4
X_14225_ _09264_ _09449_ _05012_ _05126_ _05125_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__o221ai_2
XFILLER_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11368_ _02272_ _02306_ _02307_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__nand3_4
XFILLER_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14156_ _09308_ _09406_ _04842_ _05056_ _05055_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__o221ai_4
X_13107_ _03988_ _04026_ _04028_ _04029_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nand4_1
X_10319_ term_low\[25\] term_mid\[25\] VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__nor2_1
X_11299_ _02216_ _02239_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__nand2_1
X_18964_ _09716_ _09722_ _09854_ _09855_ VGND VGND VPWR VPWR _09856_ sky130_fd_sc_hd__nand4_1
X_14087_ _04986_ _04989_ net778 net650 VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__nand4_1
X_17915_ _08619_ net137 _08772_ VGND VGND VPWR VPWR _08774_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13038_ net634 net885 VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__and2_1
X_18895_ _09781_ _09782_ _09775_ VGND VGND VPWR VPWR _09787_ sky130_fd_sc_hd__nand3_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17846_ _08663_ _08628_ VGND VGND VPWR VPWR _08707_ sky130_fd_sc_hd__nand2_1
XFILLER_67_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_93_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17777_ _08494_ _08635_ _08636_ _08634_ VGND VGND VPWR VPWR _08639_ sky130_fd_sc_hd__o211a_1
X_19516_ _00561_ _00576_ _00706_ _00705_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__a22o_4
X_14989_ _05887_ _05262_ _05260_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__nand3_4
X_16728_ _07597_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__nand2_1
X_16659_ net876 net541 _07527_ net970 VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__a22o_1
X_19447_ _00628_ _00589_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__nand2_1
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19378_ net204 _00543_ _00551_ _00553_ _00542_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__o2111ai_2
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18329_ _09045_ _09082_ VGND VGND VPWR VPWR _09179_ sky130_fd_sc_hd__nand2_1
XFILLER_147_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer229 net1025 VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_116_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap363 _02045_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_1
Xmax_cap341 _08178_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__buf_2
X_20222_ _01463_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__and2_1
Xmax_cap330 _01317_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__buf_1
Xmax_cap385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XFILLER_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap374 _08912_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_2
Xmax_cap396 _03741_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_1
X_20153_ _01389_ net215 net251 VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__a21o_1
XFILLER_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_31_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20084_ _01215_ _01232_ _01233_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__a21bo_1
XFILLER_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10670_ p_hl\[6\] p_lh\[6\] _01700_ _01705_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__o211ai_2
XFILLER_9_419 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12340_ _03268_ _03269_ _03253_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a21o_1
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12271_ _03201_ _03202_ _03203_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__and3_1
XFILLER_134_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11222_ _02078_ _02080_ _02083_ VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__o21ai_1
X_14010_ net351 _04872_ _04908_ _04910_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_147_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11153_ _02086_ _02090_ _02092_ _02072_ _02071_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_8_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11084_ net403 _02025_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__nor2_1
X_15961_ _06644_ _06726_ net173 _06836_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__o211ai_2
XFILLER_49_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15892_ _06766_ _06754_ _06765_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__nand3_2
X_17700_ net1054 net490 VGND VGND VPWR VPWR _08563_ sky130_fd_sc_hd__nand2_1
X_18680_ _09558_ _09561_ VGND VGND VPWR VPWR _09562_ sky130_fd_sc_hd__nand2_2
X_14912_ _05806_ _05808_ _05809_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__a21oi_1
XFILLER_84_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17631_ net560 net555 net500 net494 VGND VGND VPWR VPWR _08495_ sky130_fd_sc_hd__nand4_1
X_14843_ _05739_ _05737_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__nand2_4
XFILLER_90_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11986_ net324 _02878_ _02916_ _02917_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__o211a_1
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17562_ _08420_ _08414_ _08382_ _08419_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_67_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14774_ net761 net636 VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__nand2_2
X_10937_ net707 net530 net1052 net713 VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__a22oi_2
X_16513_ _07229_ _07235_ _07232_ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__a21oi_1
X_17493_ _08283_ _08355_ _08356_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_67_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13725_ net752 net694 net689 net757 VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__a22oi_4
XFILLER_17_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19301_ _10013_ _10016_ net898 net1065 _00469_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__o2111ai_4
X_16444_ _09166_ _09668_ _07313_ _07315_ VGND VGND VPWR VPWR _07317_ sky130_fd_sc_hd__or4_1
X_13656_ _04564_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__inv_2
X_19232_ net216 net717 net1128 _10125_ VGND VGND VPWR VPWR _10131_ sky130_fd_sc_hd__nand4b_1
X_10868_ net793 net1328 VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__and2_1
XFILLER_129_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12607_ net906 net995 VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19163_ _10046_ _10047_ _10039_ _10040_ VGND VGND VPWR VPWR _10056_ sky130_fd_sc_hd__o211ai_2
X_16375_ net583 net1004 net1105 net523 _07246_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__a41o_1
X_10799_ p_hl\[26\] net1306 VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__xor2_1
XFILLER_83_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18114_ _08959_ _08960_ VGND VGND VPWR VPWR _08962_ sky130_fd_sc_hd__or2_1
X_13587_ _09220_ _09417_ _04337_ _04403_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__o22a_1
XFILLER_129_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12538_ _03467_ _03338_ _03332_ VGND VGND VPWR VPWR _03470_ sky130_fd_sc_hd__nand3b_2
X_19094_ _09979_ _09981_ _09982_ VGND VGND VPWR VPWR _09985_ sky130_fd_sc_hd__and3_1
XFILLER_8_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15326_ _06195_ _06197_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__nand2_1
XFILLER_145_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18045_ _09690_ _08891_ _08894_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__and3_1
X_12469_ net679 net483 _03398_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__a21o_1
X_15257_ net726 net722 net837 a_h\[12\] VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__nand4_2
XFILLER_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14208_ _05073_ _05080_ _05108_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_111_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15188_ _05913_ _06035_ _06036_ _06005_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__a31o_1
X_14139_ net728 net724 VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__nand2_8
X_19996_ _01220_ _01221_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__nand2_1
XFILLER_101_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18947_ _09789_ _09790_ _09835_ _09837_ VGND VGND VPWR VPWR _09839_ sky130_fd_sc_hd__a22o_1
XFILLER_66_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18878_ net335 _09621_ _09766_ _09767_ VGND VGND VPWR VPWR _09770_ sky130_fd_sc_hd__nand4_4
X_17829_ _08553_ _08629_ _08633_ VGND VGND VPWR VPWR _08690_ sky130_fd_sc_hd__o21ai_1
XFILLER_55_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20771_ clknet_leaf_60_clk _00411_ VGND VGND VPWR VPWR a_h\[9\] sky130_fd_sc_hd__dfxtp_4
XFILLER_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold441 p_hh\[12\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 p_hh\[22\] VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 p_hh\[20\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 p_ll_pipe\[5\] VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap160 _07998_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_1
XFILLER_2_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold496 p_hh_pipe\[21\] VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 p_hh\[21\] VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap182 _01441_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
X_20205_ _01396_ _01398_ _01445_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__a21oi_1
Xhold485 p_ll_pipe\[31\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20136_ _09297_ _09362_ _01371_ _01372_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__a2bb2oi_1
X_20067_ _01295_ _01298_ _09308_ _09340_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11840_ net698 net487 _02773_ _02775_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__a22o_1
X_11771_ net679 net1048 net511 net508 VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_107_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ p_hl\[16\] p_lh\[16\] VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__xnor2_1
X_13510_ net777 net675 VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14490_ _05387_ _05388_ _05377_ _05378_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__o211ai_2
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ net794 _01695_ _01696_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ net1058 net785 net675 net673 VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__nand4_2
X_16160_ _07031_ net380 net1107 _06912_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__o211a_1
X_10584_ net795 net1297 VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__and2_1
X_13372_ net787 net675 VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nand2_1
X_16091_ _06966_ _06955_ _06965_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__and3_1
X_12323_ _03007_ _03149_ _03152_ _03148_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__a22o_1
Xclkload19 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_12
X_15111_ _05939_ _06007_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__nand2_1
XFILLER_126_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15042_ net723 net863 VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__nand2_1
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12254_ net682 net489 VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__nand2_1
XFILLER_5_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11205_ _02145_ _02146_ _02147_ net796 VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__a211oi_1
X_12185_ _02815_ _02816_ _02963_ _02812_ VGND VGND VPWR VPWR _03120_ sky130_fd_sc_hd__a22oi_1
X_19850_ _01057_ _01063_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__nand2_1
X_11136_ net671 net965 VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__nand2_2
X_18801_ net606 net1111 net458 _09454_ _09451_ VGND VGND VPWR VPWR _09694_ sky130_fd_sc_hd__a32o_2
X_19781_ _00877_ _00987_ _00989_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__and3_1
X_16993_ net172 _07851_ _07860_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__o21ai_2
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18732_ _09538_ _09599_ net447 _09617_ VGND VGND VPWR VPWR _09618_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15944_ _06819_ _06820_ _06749_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__a21oi_1
X_11067_ _02005_ _02008_ net967 net1106 VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__and4_1
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15875_ _06677_ _06683_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__nand2_1
X_18663_ _09533_ _09538_ _09539_ VGND VGND VPWR VPWR _09543_ sky130_fd_sc_hd__nand3_1
X_17614_ _08475_ _08477_ VGND VGND VPWR VPWR _08478_ sky130_fd_sc_hd__nand2_1
X_18594_ _09199_ _09210_ net457 _09330_ _09333_ VGND VGND VPWR VPWR _09467_ sky130_fd_sc_hd__o32a_1
XFILLER_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14826_ _05720_ _05721_ _05724_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__nand3_4
X_17545_ _08408_ _08390_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__nand2_1
XFILLER_64_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14757_ _05537_ _05656_ _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__nand3b_4
X_11969_ _02901_ _02894_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__nand2_1
X_13708_ net456 _04609_ _04607_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__o21ai_1
X_17476_ _09231_ _09679_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__nor2_1
X_14688_ _05565_ _05583_ _05564_ _05586_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__o211ai_2
X_16427_ _07295_ _07296_ _07300_ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__nand3_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13639_ _04500_ _04501_ _04502_ _04543_ net1129 VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__o2111ai_4
X_19215_ _10107_ _10106_ VGND VGND VPWR VPWR _10112_ sky130_fd_sc_hd__nand2_2
XFILLER_118_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16358_ net570 net533 net529 net572 VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__a22oi_1
XFILLER_9_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19146_ b_l\[2\] net552 net549 net1086 VGND VGND VPWR VPWR _10038_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15309_ _06086_ _06083_ _06085_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__a21bo_1
X_16289_ _07163_ _07062_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__nand2_1
XFILLER_118_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19077_ _09922_ _09923_ _09958_ _09959_ VGND VGND VPWR VPWR _09968_ sky130_fd_sc_hd__a22o_1
XFILLER_132_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18028_ _09155_ _09188_ _08873_ _08874_ VGND VGND VPWR VPWR _08878_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_93_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19979_ net568 net1043 VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_105_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20754_ clknet_leaf_49_clk _00394_ VGND VGND VPWR VPWR p_ll\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire607 net929 VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_114_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20685_ clknet_leaf_57_clk _00325_ VGND VGND VPWR VPWR p_hl\[19\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_102_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_123_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20119_ net794 _01353_ _01355_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__and3_1
X_13990_ _04893_ _04894_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__nand2_2
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12941_ _03862_ _03866_ _03868_ VGND VGND VPWR VPWR _03869_ sky130_fd_sc_hd__a21oi_1
XFILLER_58_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15660_ _06540_ _06539_ _06534_ VGND VGND VPWR VPWR _06541_ sky130_fd_sc_hd__a21oi_2
X_12872_ _03762_ _03768_ _03797_ VGND VGND VPWR VPWR _03800_ sky130_fd_sc_hd__nand3_2
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11823_ _02700_ _02756_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__nand2_2
XFILLER_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14611_ _05509_ _05510_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__and3_1
X_15591_ _06439_ _06437_ _06442_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__a21boi_1
X_17330_ _08116_ _08196_ VGND VGND VPWR VPWR _08197_ sky130_fd_sc_hd__nand2_1
XFILLER_73_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11754_ _02571_ _02691_ net796 VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_132_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14542_ net767 net642 net1135 net771 VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__a22oi_2
X_11685_ _02611_ _02616_ _02620_ _02617_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o211ai_1
X_17261_ _07962_ _08087_ _08123_ _08124_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__a2bb2oi_2
X_10705_ _01739_ _01737_ net796 VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__a21oi_1
X_14473_ _05364_ _05365_ _05325_ _05329_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__o211ai_2
X_16212_ _06847_ _07029_ net421 _07081_ _07084_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__o311ai_4
X_10636_ p_lh\[2\] p_hl\[2\] VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__and2b_1
X_17192_ _08054_ _08057_ _08051_ VGND VGND VPWR VPWR _08060_ sky130_fd_sc_hd__a21oi_2
X_13424_ _04280_ _04295_ _04293_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a21oi_2
X_19000_ _09886_ net732 net887 VGND VGND VPWR VPWR _09891_ sky130_fd_sc_hd__nand3_1
X_16143_ _07017_ _06974_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__nand2_2
XFILLER_10_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13355_ _04261_ _04262_ _04264_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__o21ai_1
X_10567_ net794 net1286 VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__and2_1
X_10498_ net1343 _01653_ _01654_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__o21a_1
X_16074_ _06746_ _06934_ _06935_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__a21oi_4
XFILLER_127_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12306_ net983 _03095_ net474 _03093_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__a31o_1
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13286_ _04198_ _04199_ _04191_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__a21o_1
XFILLER_5_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12237_ _03033_ _03167_ _03168_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__nand3_2
XFILLER_5_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15025_ _05825_ _05826_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__nand2_1
X_19902_ _01109_ _01112_ VGND VGND VPWR VPWR _01122_ sky130_fd_sc_hd__nand2_2
XFILLER_123_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19833_ _00997_ _01000_ _01043_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__nand3_1
X_12168_ _03096_ _03097_ _03090_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o21ai_1
X_11119_ _02028_ _02015_ _02017_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__a21boi_1
X_16976_ _07834_ _07841_ _07843_ _07777_ VGND VGND VPWR VPWR _07846_ sky130_fd_sc_hd__o211ai_2
X_12099_ _03030_ _03032_ _02971_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19764_ _00973_ _00712_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__nor2_4
XFILLER_1_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15927_ _06696_ _06803_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__nand2_1
Xinput6 a[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_18715_ _09534_ _09535_ _09533_ VGND VGND VPWR VPWR _09599_ sky130_fd_sc_hd__o21ai_1
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19695_ net591 net725 VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__nand2_1
XFILLER_76_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18646_ _09468_ net302 _09519_ VGND VGND VPWR VPWR _09524_ sky130_fd_sc_hd__o21ai_2
XFILLER_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15858_ _06572_ _06642_ _06565_ _06566_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__and4b_1
XFILLER_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15789_ _06664_ _06667_ _06578_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__a21boi_2
X_18577_ _09355_ _09356_ _09354_ VGND VGND VPWR VPWR _09448_ sky130_fd_sc_hd__a21oi_1
XFILLER_52_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14809_ net727 net677 VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__nand2_1
XFILLER_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17528_ _08304_ _08310_ _08307_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17459_ _08313_ _08321_ _08323_ VGND VGND VPWR VPWR _08325_ sky130_fd_sc_hd__nand3_4
X_20470_ clknet_leaf_13_clk _00110_ VGND VGND VPWR VPWR term_high\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19129_ _10017_ _10019_ net589 net1148 VGND VGND VPWR VPWR _10020_ sky130_fd_sc_hd__and4_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ clknet_leaf_4_clk _00446_ VGND VGND VPWR VPWR b_h\[12\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_46_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20737_ clknet_leaf_36_clk _00377_ VGND VGND VPWR VPWR p_ll\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire415 _08393_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_1
XFILLER_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11470_ _02409_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__inv_2
XFILLER_109_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire437 _03382_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_1
X_20668_ clknet_leaf_6_clk _00308_ VGND VGND VPWR VPWR p_hl\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10421_ _01588_ _01589_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__nor2_1
XFILLER_137_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20599_ clknet_leaf_12_clk _00239_ VGND VGND VPWR VPWR p_hh_pipe\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13140_ _04017_ _04059_ _04060_ _04062_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__nand4_1
X_10352_ _01214_ _01225_ _01236_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__o21a_1
XFILLER_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13071_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__inv_2
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12022_ _02590_ _02694_ _02956_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__o21ai_1
X_10283_ _10148_ _10169_ _00493_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16830_ _07628_ _07696_ _07697_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__nand3_1
Xclone305 net555 VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__clkbuf_16
X_16761_ net561 net516 VGND VGND VPWR VPWR _07632_ sky130_fd_sc_hd__nand2_1
Xclone316 net601 VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__clkbuf_16
Xclone338 net640 VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__clkbuf_16
X_13973_ _04733_ _04875_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nand2_1
X_15712_ net542 net595 net617 net522 VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__nand4_4
X_18500_ _09357_ _09363_ _09361_ VGND VGND VPWR VPWR _09365_ sky130_fd_sc_hd__a21oi_4
X_12924_ _03844_ _03849_ _03847_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__a21oi_1
Xclone349 b_l\[4\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__clkbuf_16
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16692_ _07452_ _07561_ _07562_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__nand3_2
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19480_ _00661_ _00662_ _00664_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__and3_1
X_15643_ _06519_ _06520_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__nand2_1
X_12855_ _03714_ _03777_ _03778_ _03712_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__a31o_1
X_18431_ _09265_ _09266_ _09289_ VGND VGND VPWR VPWR _09290_ sky130_fd_sc_hd__a21oi_4
X_15574_ _06426_ _06428_ _06456_ VGND VGND VPWR VPWR _06457_ sky130_fd_sc_hd__and3_1
X_11806_ _02610_ _02738_ net1016 net535 _02737_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__o2111ai_4
X_12786_ _03624_ _03691_ _03690_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a21boi_1
X_18362_ _09173_ _09174_ net232 _09194_ VGND VGND VPWR VPWR _09214_ sky130_fd_sc_hd__a31o_1
XFILLER_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ _02669_ _02671_ _02604_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__o21ai_1
X_17313_ net593 net585 net485 net479 VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__and4_1
X_14525_ net745 net668 _05422_ _05421_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18293_ _06681_ net805 _09134_ VGND VGND VPWR VPWR _09139_ sky130_fd_sc_hd__o21a_1
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11668_ net359 _02492_ _02512_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a21boi_4
X_17244_ _08108_ _08109_ _09253_ _09646_ VGND VGND VPWR VPWR _08112_ sky130_fd_sc_hd__o2bb2ai_1
X_14456_ _05337_ _05339_ net349 _05354_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__nand4_2
XFILLER_127_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11599_ _02532_ _02533_ _02535_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__and3_1
X_17175_ net554 net550 net1023 net516 VGND VGND VPWR VPWR _08043_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_77_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _04313_ net197 _04318_ _04315_ net796 VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__a2111oi_1
X_10619_ net794 net1218 VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__and2_1
X_14387_ _05288_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_1
X_16126_ net966 net515 _06998_ _07001_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__a22oi_1
XFILLER_115_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13338_ _04250_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__inv_2
Xmax_cap704 net705 VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__buf_8
Xmax_cap737 net738 VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__buf_8
Xmax_cap715 net716 VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__buf_6
Xmax_cap726 net727 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__buf_8
X_16057_ _06925_ _06932_ _06846_ _06933_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__o211ai_4
XFILLER_6_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap759 net760 VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_8
Xmax_cap748 net749 VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_90_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13269_ net766 net705 VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__nand2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15008_ net756 net635 VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__nand2_1
XFILLER_57_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19816_ _01014_ _01026_ _01027_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__nand3_1
XFILLER_84_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19747_ _00868_ _00951_ _00952_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__nand3_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16959_ _07825_ _07826_ VGND VGND VPWR VPWR _07829_ sky130_fd_sc_hd__nand2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19678_ _00878_ _00880_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__nand2_1
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18629_ _09501_ _09502_ _09497_ VGND VGND VPWR VPWR _09506_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_11 _00434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20522_ clknet_leaf_42_clk _00162_ VGND VGND VPWR VPWR term_low\[17\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_33 _00445_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20453_ clknet_leaf_16_clk _00093_ VGND VGND VPWR VPWR term_high\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20384_ clknet_leaf_31_clk _00024_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10970_ _01885_ _01890_ _01889_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__o21a_1
XFILLER_90_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12640_ _03395_ _03407_ _03563_ _03565_ VGND VGND VPWR VPWR _03571_ sky130_fd_sc_hd__nand4_1
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12571_ _03477_ _03462_ _03464_ VGND VGND VPWR VPWR _03502_ sky130_fd_sc_hd__o21ai_1
X_14310_ _05055_ _05201_ _05209_ _05210_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__a22oi_2
Xclkbuf_leaf_50_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11522_ _02459_ _02460_ _02449_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__nand3_2
X_15290_ net284 _06182_ _06183_ net347 VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__o2bb2ai_2
Xwire256 _07282_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
X_11453_ net698 net501 VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__and2_1
X_14241_ net392 _04997_ _04993_ _04990_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__o2bb2ai_2
X_10404_ term_mid\[36\] term_high\[36\] _01572_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__a21bo_1
XFILLER_109_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14172_ _05073_ _05074_ net316 VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__a21oi_1
X_11384_ _02323_ _02223_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__nand2_1
X_13123_ _03966_ _04009_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__a21oi_1
X_18980_ _09787_ _09788_ _09785_ VGND VGND VPWR VPWR _09871_ sky130_fd_sc_hd__a21o_1
X_10335_ _01053_ _01042_ net797 VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17931_ _08761_ _08765_ _08787_ VGND VGND VPWR VPWR _08789_ sky130_fd_sc_hd__or3b_2
XFILLER_87_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10266_ term_low\[17\] term_mid\[17\] VGND VGND VPWR VPWR _10050_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_72_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _03918_ _03728_ _03917_ _03924_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__a31o_1
X_12005_ _02789_ _02939_ _02938_ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__a21oi_2
X_17862_ _08720_ _08721_ VGND VGND VPWR VPWR _08722_ sky130_fd_sc_hd__nor2_1
XFILLER_79_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16813_ _07678_ _07681_ _07682_ _07496_ VGND VGND VPWR VPWR _07684_ sky130_fd_sc_hd__o2bb2a_1
X_19601_ net835 net574 net1033 net579 VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__a22oi_2
X_10197_ net728 VGND VGND VPWR VPWR _09329_ sky130_fd_sc_hd__inv_2
XFILLER_120_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17793_ _08652_ _08653_ a_l\[10\] net472 VGND VGND VPWR VPWR _08655_ sky130_fd_sc_hd__nand4_1
X_16744_ _07610_ _07611_ _07600_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__nand3_1
Xclone168 net1115 VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__clkbuf_16
XFILLER_93_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone179 net996 VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__clkbuf_16
XFILLER_47_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19532_ _00589_ _00629_ _00723_ _00628_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__o211ai_2
X_13956_ _04858_ _04859_ _04861_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__and3_1
X_16675_ _07540_ _07541_ _07510_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__nand3_4
X_12907_ _03833_ _03834_ _03821_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__a21oi_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13887_ _04788_ _04791_ _04792_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__a21bo_1
X_19463_ net755 net567 VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__nand2_1
X_15626_ net631 net512 _06506_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__a21o_1
X_12838_ _03634_ _03651_ _03653_ _03762_ net267 VGND VGND VPWR VPWR _03767_ sky130_fd_sc_hd__o2111ai_1
X_18414_ net798 net754 VGND VGND VPWR VPWR _09271_ sky130_fd_sc_hd__nand2_1
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19394_ _00572_ _00574_ _00575_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__o21a_1
X_15557_ net528 net532 VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__nand2_8
X_12769_ _03696_ _03697_ _03612_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__nand3_1
X_18345_ _09186_ _09194_ VGND VGND VPWR VPWR _09196_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_41_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18276_ _09115_ _09120_ _09121_ VGND VGND VPWR VPWR _09122_ sky130_fd_sc_hd__nand3_2
X_14508_ _05263_ _05409_ _05410_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__o21a_1
X_15488_ _06375_ _06376_ _06368_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput31 a[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
X_17227_ net593 net485 net479 net600 VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__a22oi_2
Xinput20 a[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_14439_ _05203_ _05208_ _05205_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__a21oi_1
Xmax_cap512 net513 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_12
Xmax_cap501 b_h\[8\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_6
Xinput53 b[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 b[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput64 b[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
X_17158_ _07730_ _07881_ _07879_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__a21boi_2
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap545 net547 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__buf_12
Xmax_cap523 net524 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_114_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16109_ net586 net582 VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__nand2_8
X_17089_ _07954_ _07955_ _09242_ _09646_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__o2bb2a_1
Xmax_cap556 net557 VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__buf_12
Xmax_cap567 net568 VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__buf_12
XFILLER_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap589 net941 VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_8
XFILLER_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xload_slew795 _09690_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__buf_12
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20505_ clknet_leaf_35_clk _00145_ VGND VGND VPWR VPWR term_low\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20436_ clknet_leaf_13_clk _00076_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfxtp_1
X_20367_ clknet_leaf_47_clk _00007_ VGND VGND VPWR VPWR b_l\[7\] sky130_fd_sc_hd__dfxtp_4
XFILLER_106_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20298_ _09373_ _09384_ _01530_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__o21a_1
XFILLER_0_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ _05686_ _05687_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__nand2_1
X_13810_ _09264_ _09417_ _04715_ _04716_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__o211ai_2
X_10953_ _01875_ _01879_ _01898_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__nand4_1
X_13741_ _04644_ _04646_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__nand2_1
XFILLER_28_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ _07194_ _07198_ _07328_ _07329_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__a22o_1
XFILLER_73_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10884_ net794 net1268 VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__and2_1
X_13672_ _04577_ _04576_ _04478_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__a21o_1
X_16391_ _07260_ net505 a_l\[6\] VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_23_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_12623_ _03552_ net475 net682 _03551_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__nand4_1
X_15411_ _06217_ _06303_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__nand2_1
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12554_ net176 _03485_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__nor2_2
X_18130_ net459 _06681_ _08916_ _08919_ VGND VGND VPWR VPWR _08978_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_42_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15342_ _06225_ _06226_ _06233_ _06234_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__nand4_2
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11505_ net151 _02443_ _02444_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__o21a_1
X_18061_ net627 net764 _08908_ _08909_ VGND VGND VPWR VPWR _08910_ sky130_fd_sc_hd__a22oi_4
X_15273_ _06091_ _06162_ net730 net643 _06166_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__o2111ai_2
X_17012_ _07874_ _07880_ _07879_ VGND VGND VPWR VPWR _07882_ sky130_fd_sc_hd__o21ai_1
X_12485_ net356 _03322_ _03411_ _03412_ _03321_ VGND VGND VPWR VPWR _03417_ sky130_fd_sc_hd__o2111ai_2
X_14224_ net756 net750 net670 net667 VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__nand4_1
X_11436_ _02292_ _02374_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__nand2_1
X_11367_ _02176_ _02179_ _02305_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__a21oi_1
X_14155_ _04842_ _05056_ net731 net699 _05055_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__o2111ai_1
XFILLER_98_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13106_ _03988_ _04026_ _04028_ _04029_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__and4_1
X_18963_ _09852_ _09853_ _09739_ VGND VGND VPWR VPWR _09855_ sky130_fd_sc_hd__a21bo_1
X_14086_ net778 net650 _04986_ _04989_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__a22o_1
X_10318_ net794 _00849_ _00870_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__and3_1
XFILLER_140_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11298_ _02151_ _02217_ _02218_ _02224_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__a31o_1
X_17914_ _08619_ net137 _08772_ VGND VGND VPWR VPWR _08773_ sky130_fd_sc_hd__o21a_1
X_13037_ _03961_ net478 net839 _03960_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__nand4_4
X_10249_ _09690_ net1245 VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__and2_1
XFILLER_67_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18894_ _09644_ _09774_ _09783_ _09784_ VGND VGND VPWR VPWR _09786_ sky130_fd_sc_hd__o211ai_2
XFILLER_93_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17845_ _08704_ _08705_ VGND VGND VPWR VPWR _08706_ sky130_fd_sc_hd__nand2_1
XFILLER_39_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17776_ _08566_ _08563_ _08564_ _08637_ VGND VGND VPWR VPWR _08638_ sky130_fd_sc_hd__o211ai_4
X_16727_ _07593_ _07595_ _07596_ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_85_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19515_ _00701_ net230 _00702_ _00704_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__nand4_4
X_14988_ _05662_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__nor2_4
XFILLER_90_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13939_ net742 net735 net699 net695 VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__nand4_2
X_16658_ _07527_ net970 _07523_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__a21oi_2
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19446_ _00628_ _00630_ _00589_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__a21o_4
X_16589_ net812 net1032 _07459_ _07460_ VGND VGND VPWR VPWR _07461_ sky130_fd_sc_hd__a22o_1
X_15609_ _06470_ _06471_ _06489_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__nand4_1
X_19377_ net204 _00543_ _00555_ _00542_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__o211ai_2
XFILLER_34_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
X_18328_ _09172_ _09131_ VGND VGND VPWR VPWR _09178_ sky130_fd_sc_hd__nand2_1
XFILLER_147_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer208 net1053 VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_20_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18259_ _08856_ _08890_ _08950_ _09018_ VGND VGND VPWR VPWR _09106_ sky130_fd_sc_hd__or4b_1
XFILLER_147_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap342 _08114_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_4
Xmax_cap353 _03515_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_1
X_20221_ _01461_ _01462_ _09340_ _09362_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20152_ _01389_ net215 _01381_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__a21oi_1
XFILLER_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20083_ _01226_ _01227_ _01231_ _01213_ _01212_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__a311oi_2
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12270_ _03045_ _03046_ _03060_ _03062_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__o31ai_1
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20419_ clknet_leaf_27_clk _00059_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfxtp_1
X_11221_ _02161_ _02162_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__nor2_2
XFILLER_107_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11152_ _02074_ _02091_ _02092_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__and3_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ _02022_ _02023_ _02019_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__a21oi_1
X_15960_ _06644_ _06726_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15891_ _06682_ _06752_ _06763_ _06764_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__o211ai_4
XFILLER_76_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14911_ _05683_ net655 net745 _05684_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__a31oi_2
XFILLER_124_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17630_ net555 net494 VGND VGND VPWR VPWR _08494_ sky130_fd_sc_hd__nand2_4
X_14842_ _05733_ _05735_ _05736_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__a21oi_2
X_11985_ net324 _02878_ _02916_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__o21ai_2
XFILLER_91_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17561_ _08423_ _08383_ _08422_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__nand3_1
XFILLER_16_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14773_ net761 net636 VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__and2_1
X_19300_ _10013_ _10016_ _10019_ _00467_ _00469_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__o2111a_1
X_10936_ net707 net1052 _01866_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__and3_1
X_16512_ _07229_ _07235_ _07232_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__a21o_1
X_17492_ _08354_ _08350_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_67_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13724_ net757 net689 VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__nand2_1
X_10867_ net793 net1285 VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__and2_1
X_16443_ _02589_ _06441_ a_l\[0\] net477 _07314_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__o2111a_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13655_ _04558_ _04559_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__xnor2_1
X_19231_ _10121_ _10124_ net216 VGND VGND VPWR VPWR _10130_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_80_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12606_ net659 net495 VGND VGND VPWR VPWR _03537_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19162_ _10039_ _10040_ _10046_ _10047_ VGND VGND VPWR VPWR _10055_ sky130_fd_sc_hd__o2bb2ai_2
X_16374_ net586 net515 _07243_ _07245_ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__a22o_1
X_10798_ _01818_ _01819_ _01820_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__o21a_1
X_18113_ _08959_ _08960_ VGND VGND VPWR VPWR _08961_ sky130_fd_sc_hd__nor2_1
X_13586_ _09264_ _09395_ _04493_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__o211ai_2
XFILLER_12_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12537_ _03301_ _03304_ _03331_ _03468_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__o211ai_2
X_19093_ _09166_ _09384_ _09978_ _09980_ VGND VGND VPWR VPWR _09984_ sky130_fd_sc_hd__o22ai_1
X_15325_ _06211_ _06218_ _06219_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__o21a_1
XFILLER_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18044_ _08853_ _08856_ _08890_ VGND VGND VPWR VPWR _08894_ sky130_fd_sc_hd__a21o_1
X_12468_ _03398_ _03399_ VGND VGND VPWR VPWR _03400_ sky130_fd_sc_hd__nand2_1
X_15256_ net726 net722 net837 net870 VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__and4_1
XFILLER_144_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11419_ net652 net546 VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__nand2_1
X_14207_ _05073_ _05080_ _05108_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__and3_1
X_15187_ _09384_ _09460_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__nor2_1
XFILLER_141_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12399_ _03325_ _03326_ _03329_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__nand3_4
X_14138_ net728 net724 VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__and2_4
XFILLER_113_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_747 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19995_ net735 net557 net551 net742 VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__a22oi_2
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_18946_ _09828_ _09834_ _09832_ _09836_ _09793_ VGND VGND VPWR VPWR _09838_ sky130_fd_sc_hd__o221ai_2
X_14069_ net767 net662 net656 net771 VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__a22oi_4
X_18877_ _09621_ net335 _09766_ _09767_ VGND VGND VPWR VPWR _09769_ sky130_fd_sc_hd__a22o_4
XFILLER_94_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17828_ _09340_ _09657_ _08553_ _08633_ VGND VGND VPWR VPWR _08689_ sky130_fd_sc_hd__o31a_1
XFILLER_55_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17759_ _08274_ _08027_ _08619_ VGND VGND VPWR VPWR _08622_ sky130_fd_sc_hd__a21oi_2
XFILLER_81_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20770_ clknet_leaf_60_clk _00410_ VGND VGND VPWR VPWR a_h\[8\] sky130_fd_sc_hd__dfxtp_4
X_19429_ net598 net729 VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__nand2_1
XFILLER_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_136_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold420 p_ll_pipe\[23\] VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap161 _07168_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_6
XFILLER_132_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold442 p_ll\[3\] VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 term_low\[12\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 p_ll_pipe\[16\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
X_20204_ _01396_ _01398_ _01444_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__a21bo_1
Xhold464 p_hh\[9\] VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap172 _07849_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xhold475 mid_sum\[3\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 mid_sum\[10\] VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap183 _00693_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_2
Xmax_cap194 _05240_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_129_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold497 p_ll\[13\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20135_ _01283_ _01369_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__nand2_2
XFILLER_98_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20066_ _01218_ _01296_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__nand2_1
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net672 net508 VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__nand2_2
XFILLER_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10721_ _01751_ _01752_ _01753_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__o21a_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13440_ _04287_ _04349_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__nand2_2
X_10652_ _01691_ _01692_ _01694_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ net793 net1255 VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__and2_1
XFILLER_139_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13371_ net777 net986 VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__nand2_1
X_16090_ _06960_ _06962_ _06957_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ _03007_ _03149_ _03152_ _03148_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a22oi_2
X_15110_ net726 net663 VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__nand2_1
X_12253_ net679 net672 net499 net492 VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__nand4_2
X_15041_ net723 net956 VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__nand2_1
X_11204_ _02060_ _02138_ _02142_ _02146_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__a31oi_4
XFILLER_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12184_ _02817_ _02818_ _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__nand3_1
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16992_ _07849_ _07851_ _07860_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__o21bai_1
X_11135_ net681 net534 VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__nand2_1
XFILLER_68_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18800_ _09688_ _09692_ VGND VGND VPWR VPWR _09693_ sky130_fd_sc_hd__nand2_1
X_19780_ net366 _00987_ _00990_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__a21oi_1
X_15943_ _06709_ _06712_ _06818_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__nand3_2
X_11066_ _09428_ _09592_ _02009_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__o21ai_1
X_18731_ _04555_ _06521_ _09609_ VGND VGND VPWR VPWR _09617_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15874_ _06678_ _06679_ _06677_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__a21oi_2
X_18662_ _09538_ _09539_ _09533_ VGND VGND VPWR VPWR _09542_ sky130_fd_sc_hd__a21o_1
XFILLER_49_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17613_ _08470_ _08471_ net941 net472 VGND VGND VPWR VPWR _08477_ sky130_fd_sc_hd__nand4_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18593_ net610 net604 net458 net1148 net619 VGND VGND VPWR VPWR _09466_ sky130_fd_sc_hd__a32o_1
X_14825_ _05613_ _05614_ _05617_ _05612_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__a22oi_2
X_17544_ _08391_ _08405_ _08407_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__nand3_1
X_14756_ net163 _05652_ _05538_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__a21o_1
X_11968_ _02895_ _02900_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__nand2_2
X_13707_ _09220_ _09439_ net456 _04609_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__o22a_1
X_10919_ net1062 _01860_ _01859_ _01861_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__o22ai_1
X_11899_ _02774_ _02833_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__nand2_2
X_17475_ _08230_ _08235_ _08337_ _08338_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__and4_1
X_19214_ _10074_ _10104_ _10106_ VGND VGND VPWR VPWR _10111_ sky130_fd_sc_hd__and3_1
X_14687_ _05566_ _05581_ _05583_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__nand3_1
X_16426_ net281 _07166_ _07165_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__a21boi_1
X_13638_ _04544_ _04543_ _04503_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a21o_1
X_16357_ net570 net533 VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__nand2_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13569_ _04477_ _04478_ _04389_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__a21oi_4
X_19145_ b_l\[2\] net552 net549 net1086 VGND VGND VPWR VPWR _10037_ sky130_fd_sc_hd__a22oi_2
XFILLER_117_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19076_ _09922_ _09923_ _09958_ _09959_ VGND VGND VPWR VPWR _09967_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_30_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15308_ _06130_ _06135_ _06199_ _06200_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__a22o_1
XFILLER_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16288_ _07156_ _07155_ _07088_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__a21o_1
X_18027_ _08873_ _08874_ _08869_ VGND VGND VPWR VPWR _08877_ sky130_fd_sc_hd__a21o_1
XFILLER_126_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15239_ _06089_ _06131_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__nand2_2
XFILLER_99_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19978_ net580 net721 VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__nand2_1
X_18929_ _09155_ _09319_ _09658_ _09816_ _09815_ VGND VGND VPWR VPWR _09821_ sky130_fd_sc_hd__o221ai_2
XFILLER_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20753_ clknet_leaf_49_clk _00393_ VGND VGND VPWR VPWR p_ll\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ clknet_leaf_57_clk _00324_ VGND VGND VPWR VPWR p_hl\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20118_ _01345_ _01350_ _01351_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__nand3b_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12940_ net680 _03720_ net474 _03718_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__a31o_1
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20049_ _01200_ _01255_ _01254_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__o21a_1
X_12871_ _03736_ _03739_ _03763_ _03798_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__o211ai_4
X_11822_ _02758_ _02699_ _02757_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__nand3_4
X_14610_ _01888_ net455 net390 _05362_ _05369_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__o2111ai_4
X_15590_ _06470_ _06471_ VGND VGND VPWR VPWR _06472_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_64_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11753_ _02689_ _02690_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__nand2_1
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14541_ net767 net642 VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__nand2_1
X_11684_ _02618_ _02619_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__a21oi_1
X_17260_ _08125_ _08124_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__nand2_1
X_10704_ p_hl\[11\] p_lh\[11\] _01737_ _01738_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__o211ai_1
X_14472_ _05325_ _05329_ _05366_ _05370_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__o2bb2ai_2
X_16211_ _07081_ _07084_ _07032_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__a21bo_2
X_10635_ p_hl\[2\] p_lh\[2\] VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__and2b_1
X_17191_ _08054_ _08057_ _09297_ _09613_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__o2bb2ai_1
X_13423_ _04294_ _04299_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__nand2_1
X_16142_ _06972_ _06973_ _07014_ _07016_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__nand4_2
X_13354_ net714 net963 net1125 _04262_ _04264_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__a311o_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ _03236_ _03235_ _03234_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__nand3_2
XFILLER_6_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10566_ net794 net1289 VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__and2_1
X_10497_ _01653_ net1343 net796 VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__a21oi_1
X_16073_ _06937_ _06938_ _06832_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__a21oi_2
X_13285_ _04162_ _04195_ net777 net700 _04194_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__o2111ai_2
X_12236_ net293 _03028_ _03165_ _03166_ VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__a22oi_4
XFILLER_5_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19901_ net332 VGND VGND VPWR VPWR _01121_ sky130_fd_sc_hd__inv_2
X_15024_ _05810_ _05807_ _05806_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__o21ai_2
X_12167_ net177 _03089_ net199 _03088_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_75_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19832_ _00997_ _01041_ _01043_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__nand3_1
X_11118_ _02028_ _02015_ _02011_ _02016_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16975_ _07834_ _07841_ _07843_ _07777_ VGND VGND VPWR VPWR _07845_ sky130_fd_sc_hd__o211a_1
X_12098_ net293 _03028_ VGND VGND VPWR VPWR _03033_ sky130_fd_sc_hd__nand2_1
XFILLER_68_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19763_ _00707_ _00708_ _00853_ _00854_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__nand4_4
X_11049_ _01993_ _01992_ _01990_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__a21o_1
X_15926_ _06692_ _06695_ _06697_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__o21ai_2
Xinput7 a[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18714_ _05043_ net847 _09597_ VGND VGND VPWR VPWR _09598_ sky130_fd_sc_hd__a21oi_2
X_19694_ _00750_ _00759_ _00763_ _00757_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15857_ _06734_ _06735_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__nand2_1
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18645_ _09519_ _09473_ VGND VGND VPWR VPWR _09523_ sky130_fd_sc_hd__nand2_2
XFILLER_92_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14808_ _05706_ _05707_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__nand2_1
X_15788_ _06656_ _06665_ _06666_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__nand3_2
X_18576_ net922 _06867_ _09354_ VGND VGND VPWR VPWR _09447_ sky130_fd_sc_hd__o21ai_1
X_17527_ _08304_ _08310_ _08307_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__a21o_1
X_14739_ _05596_ _05598_ _05636_ _05638_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__nand4_4
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17458_ net340 _08317_ _08320_ _08322_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_TAPCELL_ROW_15_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16409_ _07256_ _07257_ _07279_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__nand3_1
X_17389_ _08250_ _08251_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__nand2_1
X_19128_ net579 net755 net760 net575 VGND VGND VPWR VPWR _10019_ sky130_fd_sc_hd__nand4_4
X_19059_ _09937_ _09938_ _09947_ _09948_ VGND VGND VPWR VPWR _09950_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_102_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20805_ clknet_leaf_4_clk _00445_ VGND VGND VPWR VPWR b_h\[11\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_46_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20736_ clknet_leaf_32_clk _00376_ VGND VGND VPWR VPWR p_ll\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ term_mid\[40\] term_high\[40\] VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_137_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20667_ clknet_leaf_24_clk _00307_ VGND VGND VPWR VPWR p_hl\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire427 _05558_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_1
X_20598_ clknet_leaf_13_clk _00238_ VGND VGND VPWR VPWR p_hh_pipe\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10351_ _01225_ _01214_ net797 VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__a21oi_1
X_13070_ _03994_ _03995_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__nand2_1
X_10282_ _00471_ _00482_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__nand2_1
X_12021_ _02955_ _02695_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__nand2_1
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16760_ _07519_ _07538_ _07536_ _07530_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o2bb2ai_4
X_13972_ net1122 net667 net660 net771 VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a22oi_2
X_15711_ _06588_ _06589_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__nand2_2
X_12923_ _03849_ _03844_ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__nand2_1
X_16691_ _07452_ _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__nand2_1
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18430_ _09285_ _09288_ VGND VGND VPWR VPWR _09289_ sky130_fd_sc_hd__nand2_4
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15642_ net1083 net531 net527 net1120 VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__a22oi_4
X_12854_ _03714_ _03777_ _03778_ VGND VGND VPWR VPWR _03783_ sky130_fd_sc_hd__nand3_1
X_15573_ _06454_ _06455_ VGND VGND VPWR VPWR _06456_ sky130_fd_sc_hd__nand2_1
X_11805_ _02737_ _02739_ _09504_ _09592_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_92_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12785_ _03690_ _03713_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__nand2_1
X_18361_ _09173_ _09174_ net232 _09194_ VGND VGND VPWR VPWR _09213_ sky130_fd_sc_hd__a31oi_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11736_ _02669_ _02671_ _02604_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__o21bai_4
X_17312_ _08178_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__inv_2
X_18292_ _09050_ _09135_ VGND VGND VPWR VPWR _09138_ sky130_fd_sc_hd__nand2_1
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14524_ _05421_ _05422_ net745 net668 VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_32_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _08108_ _08109_ _08104_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__a21o_1
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11667_ _02492_ net997 _02506_ _02511_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__o2bb2ai_4
X_14455_ _05340_ _05354_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__nand2_1
XFILLER_128_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11598_ _02532_ _02533_ _02534_ _02398_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__o2bb2ai_1
X_17174_ net554 net550 net1023 net516 VGND VGND VPWR VPWR _08042_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_77_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _04255_ _04209_ _04178_ _04312_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__nor4b_4
X_10618_ net794 net1176 VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__and2_1
X_14386_ _05161_ _05166_ _05284_ _05286_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nand4_4
X_10549_ net793 net1290 VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__and2_1
XFILLER_128_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16125_ net595 net570 net1063 net521 VGND VGND VPWR VPWR _07001_ sky130_fd_sc_hd__nand4_2
X_13337_ _04248_ _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__nand2_1
Xmax_cap705 a_h\[2\] VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__buf_8
XFILLER_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap716 b_l\[15\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__buf_8
Xmax_cap727 net728 VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__buf_12
XFILLER_143_758 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16056_ _06926_ _06927_ net238 VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__a21o_1
Xmax_cap738 b_l\[10\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_8
Xmax_cap749 b_l\[8\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_90_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13268_ net772 net953 VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__nand2_8
X_15007_ net745 _05796_ net649 _05798_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__a31o_1
XFILLER_111_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12219_ _09504_ _09602_ _03008_ _03151_ _03150_ VGND VGND VPWR VPWR _03153_ sky130_fd_sc_hd__o221ai_2
X_13199_ _04118_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19815_ _01024_ _01025_ _01013_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__a21oi_2
X_16958_ _07652_ _07816_ _07824_ _07815_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__o211ai_2
X_19746_ _00949_ _00950_ _00869_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__a21oi_4
X_15909_ _06786_ _06785_ _06750_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__nand3_4
XFILLER_37_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16889_ _07755_ net488 net600 VGND VGND VPWR VPWR _07759_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_88_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19677_ _00877_ net1013 net893 _00875_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__nand4_2
XFILLER_92_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18628_ _09501_ _09502_ _09498_ VGND VGND VPWR VPWR _09505_ sky130_fd_sc_hd__a21oi_1
X_18559_ _09424_ _09425_ _09323_ VGND VGND VPWR VPWR _09430_ sky130_fd_sc_hd__nand3_2
XFILLER_80_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 _00435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20521_ clknet_leaf_42_clk _00161_ VGND VGND VPWR VPWR term_low\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_23 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_34 net713 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20452_ clknet_leaf_16_clk _00092_ VGND VGND VPWR VPWR term_high\[44\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20383_ clknet_leaf_31_clk _00023_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12570_ _03463_ _03476_ _03464_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a21boi_2
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11521_ _01871_ _02338_ net708 net487 _02456_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__o2111ai_1
X_20719_ clknet_leaf_23_clk _00359_ VGND VGND VPWR VPWR p_lh\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire257 _07224_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_2
X_11452_ _02296_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__nand2_1
Xwire246 _03417_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14240_ net315 _05141_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__nor2_1
X_10403_ _01573_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__nor2_1
X_11383_ _02322_ _02323_ _02220_ _02221_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_59_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14171_ _04854_ _04838_ _04849_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__a21boi_1
X_13122_ _04044_ _04045_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__nand2_1
X_10334_ term_low\[26\] net1370 _01021_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__a21bo_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17930_ _08761_ _08765_ _08787_ VGND VGND VPWR VPWR _08788_ sky130_fd_sc_hd__o21ba_1
XFILLER_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10265_ term_low\[16\] net1316 _10029_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_72_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _03918_ _03728_ _03917_ _03924_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__a31oi_1
X_12004_ _02764_ _02767_ _02789_ _02939_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__o211a_1
X_17861_ _08718_ _08719_ _09340_ _09668_ VGND VGND VPWR VPWR _08721_ sky130_fd_sc_hd__o2bb2a_1
X_10196_ net564 VGND VGND VPWR VPWR _09319_ sky130_fd_sc_hd__inv_8
XFILLER_120_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16812_ _07494_ _07499_ _07496_ VGND VGND VPWR VPWR _07683_ sky130_fd_sc_hd__a21oi_2
X_19600_ net835 net574 VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__nand2_1
X_17792_ _08652_ _08653_ VGND VGND VPWR VPWR _08654_ sky130_fd_sc_hd__nand2_1
Xclone125 net772 net1020 VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__nand2_4
Xclone147 net959 VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__clkbuf_16
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19531_ _00610_ _00614_ _00615_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__a21oi_1
X_16743_ _07601_ _07612_ _07613_ VGND VGND VPWR VPWR _07614_ sky130_fd_sc_hd__nand3_2
Xclone169 net988 VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__clkbuf_16
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13955_ _04719_ _04725_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__nand2_1
X_16674_ _07511_ _07542_ _07543_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__nand3_2
X_12906_ _09635_ _03826_ net884 net976 _03829_ VGND VGND VPWR VPWR _03834_ sky130_fd_sc_hd__o2111ai_2
X_13886_ _09177_ _09329_ _04788_ _04791_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o211ai_1
X_19462_ net878 net562 VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__nand2_1
X_15625_ net631 _06466_ net515 _06468_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__a31o_1
X_12837_ _03762_ net267 _03764_ _03654_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__o2bb2ai_1
X_18413_ net1100 net1148 VGND VGND VPWR VPWR _09270_ sky130_fd_sc_hd__nand2_1
XFILLER_61_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19393_ _00572_ _00574_ net797 VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__a21oi_1
X_18344_ _09191_ _09193_ VGND VGND VPWR VPWR _09195_ sky130_fd_sc_hd__nand2_1
X_15556_ _06413_ _06438_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__nand2_2
X_12768_ _03696_ _03697_ _03612_ VGND VGND VPWR VPWR _03698_ sky130_fd_sc_hd__a21o_1
XFILLER_61_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11719_ _02484_ _02489_ _02655_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__a22oi_4
X_12699_ _03625_ _03626_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__nand2_1
X_18275_ _09117_ net754 net1100 VGND VGND VPWR VPWR _09121_ sky130_fd_sc_hd__nand3_1
X_14507_ _05263_ _05409_ net65 VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__a21oi_1
X_15487_ _06352_ _06353_ _06375_ _06376_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__o22a_1
X_17226_ net606 net476 VGND VGND VPWR VPWR _08094_ sky130_fd_sc_hd__nand2_1
Xinput10 a[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput21 a[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
X_14438_ _05203_ _05208_ _05205_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__a21o_1
XFILLER_30_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 a[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
X_17157_ _07874_ _07880_ _07730_ VGND VGND VPWR VPWR _08026_ sky130_fd_sc_hd__o21ai_1
Xmax_cap502 net503 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__buf_8
Xinput54 b[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput43 b[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap535 net536 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__buf_8
Xmax_cap513 net514 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_6
Xmax_cap524 b_h\[4\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_12
Xinput65 rst VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_16
X_14369_ net767 net649 VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__nand2_1
X_16108_ _09253_ _09275_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap546 net547 VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__buf_8
X_17088_ _07954_ _07955_ _07952_ VGND VGND VPWR VPWR _07957_ sky130_fd_sc_hd__a21o_1
Xmax_cap557 net560 VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__buf_8
Xmax_cap579 net580 VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__buf_12
X_16039_ _06858_ _06888_ _06889_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__nand3_4
XFILLER_124_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19729_ _00909_ _00910_ _00931_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__o21ai_4
XFILLER_92_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20504_ clknet_leaf_15_clk _00144_ VGND VGND VPWR VPWR term_mid\[48\] sky130_fd_sc_hd__dfxtp_1
XFILLER_147_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20435_ clknet_leaf_14_clk _00075_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfxtp_1
XFILLER_106_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20366_ clknet_leaf_49_clk _00006_ VGND VGND VPWR VPWR b_l\[6\] sky130_fd_sc_hd__dfxtp_4
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20297_ _01542_ _01521_ net794 _01543_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_54_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10952_ _01883_ _01884_ _01896_ _01897_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__o211ai_1
XFILLER_56_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13740_ _04627_ net393 _04642_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__and3_1
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ _04579_ _04578_ _04382_ _04476_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__o2bb2ai_2
X_10883_ net794 net1236 VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__and2_1
X_15410_ _06214_ _06215_ _06302_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__a21boi_1
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16390_ _07131_ net513 a_l\[7\] VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__nand3_1
X_12622_ net684 net475 VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__nand2_1
XFILLER_73_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12553_ _03346_ _03480_ _03481_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__nand3_4
X_15341_ _06225_ _06226_ _06233_ _06234_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11504_ _02442_ _02443_ net796 VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__a21oi_1
X_18060_ net623 net615 net774 net769 VGND VGND VPWR VPWR _08909_ sky130_fd_sc_hd__nand4_4
X_15272_ _06091_ _06162_ _06160_ _06166_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__o211a_1
X_17011_ _07719_ _07877_ _07876_ _07875_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__o211ai_2
X_12484_ _03411_ _03414_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__nand2_1
X_14223_ net756 net750 net670 net667 VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__and4_1
X_11435_ net1048 net525 net1059 net1061 VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__a22oi_1
X_11366_ _02288_ _02289_ _02298_ _02300_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__nand4_2
X_14154_ _05055_ _05058_ _09308_ _09406_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__o2bb2ai_1
X_11297_ _02148_ _02237_ _02238_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__o21a_1
XFILLER_98_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13105_ _04026_ _04028_ _04029_ _03988_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__a22o_1
X_18962_ _09736_ _09738_ net987 _09850_ _09852_ VGND VGND VPWR VPWR _09854_ sky130_fd_sc_hd__o221ai_4
X_14085_ net778 net650 _04986_ _04989_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__a22oi_4
X_10317_ term_low\[23\] term_mid\[23\] _00827_ _00838_ VGND VGND VPWR VPWR _00870_
+ sky130_fd_sc_hd__o211ai_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10248_ _09690_ net1189 VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__and2_1
X_17913_ _08614_ _08669_ _08771_ VGND VGND VPWR VPWR _08772_ sky130_fd_sc_hd__and3_1
X_13036_ _03960_ _03961_ _09493_ _09668_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__o2bb2ai_1
X_18893_ _09781_ _09782_ _09775_ VGND VGND VPWR VPWR _09785_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17844_ _08647_ _08651_ _08653_ _08701_ _08702_ VGND VGND VPWR VPWR _08705_ sky130_fd_sc_hd__o2111ai_1
XFILLER_66_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17775_ _08494_ _08635_ _08636_ VGND VGND VPWR VPWR _08637_ sky130_fd_sc_hd__o21ai_1
X_14987_ _05775_ _05659_ _05658_ _05777_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__nand4_4
X_16726_ _09144_ _09668_ _07593_ _07595_ VGND VGND VPWR VPWR _07597_ sky130_fd_sc_hd__o211ai_2
XFILLER_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19514_ _00701_ _00702_ _00703_ _00549_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__o2bb2ai_4
X_13938_ _04841_ _04842_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__nand2_1
XFILLER_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19445_ _00626_ _00627_ _00591_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__nand3_4
X_16657_ _07527_ net970 VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__nand2_1
X_13869_ _04770_ _04765_ _04653_ _04771_ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__o211ai_4
X_16588_ net928 a_l\[6\] net496 net491 VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__nand4_2
X_15608_ _06485_ _06487_ _06473_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__nand3_4
X_19376_ _00542_ _00544_ _00555_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__a21o_1
X_15539_ _09188_ _09526_ _06421_ _06422_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__o211ai_2
X_18327_ _09126_ _09127_ _09170_ net1089 VGND VGND VPWR VPWR _09176_ sky130_fd_sc_hd__o211ai_2
XFILLER_147_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer209 net1005 VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd1_1
X_18258_ net219 _09018_ _09097_ _09103_ VGND VGND VPWR VPWR _09105_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_20_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17209_ _08049_ _07907_ _08048_ _08075_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__o211ai_4
XFILLER_128_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18189_ _09030_ _09033_ _09035_ VGND VGND VPWR VPWR _09036_ sky130_fd_sc_hd__a21oi_1
Xmax_cap310 _05914_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_1
XFILLER_116_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap343 _07935_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
X_20220_ _01461_ _01462_ net557 b_l\[14\] VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__nand4_1
Xmax_cap332 _01120_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__buf_6
XFILLER_131_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap387 _06581_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_6
Xmax_cap376 _07793_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_1
X_20151_ _01387_ _01388_ _09286_ _09384_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_85_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20082_ _01312_ _01313_ _01101_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__nand3_2
XFILLER_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20418_ clknet_leaf_18_clk _00058_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11220_ _02064_ _02159_ _02154_ _02158_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__o211a_4
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11151_ _02093_ _02073_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__nand2_1
X_20349_ net794 net46 VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__and2_1
XFILLER_1_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _02019_ _02022_ _02023_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__and3_1
XFILLER_103_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15890_ _06682_ _06752_ _06763_ _06764_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__o211a_1
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14910_ net745 _05683_ net655 _05684_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__a31o_1
XFILLER_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14841_ _05621_ _05626_ _05728_ _05734_ _05733_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__o221ai_4
X_17560_ _08419_ _08421_ _08382_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__a21oi_2
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11984_ _02919_ _02880_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__nand2_1
X_16511_ _07379_ _07371_ VGND VGND VPWR VPWR _07384_ sky130_fd_sc_hd__nand2_1
X_14772_ net312 _05587_ _05588_ _05562_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__a31oi_4
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10935_ net795 _01881_ _01882_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__and3_1
X_17491_ _08285_ _08339_ _08348_ _08349_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_71_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13723_ net748 net701 VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__nand2_1
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10866_ net793 net1305 VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__and2_1
X_16442_ a_l\[2\] net628 net484 net480 VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__and4_1
X_13654_ net714 net963 _04554_ _04557_ _04560_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__a311o_1
X_19230_ _10124_ net216 _10121_ VGND VGND VPWR VPWR _10129_ sky130_fd_sc_hd__o21ai_1
X_16373_ net587 net515 _07243_ _07245_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_80_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12605_ net920 net489 VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__nand2_1
X_19161_ _10053_ _10040_ _10039_ VGND VGND VPWR VPWR _10054_ sky130_fd_sc_hd__nand3_1
X_10797_ _01819_ _01818_ net796 VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__a21oi_1
X_18112_ _08957_ _08958_ VGND VGND VPWR VPWR _08960_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15324_ _06218_ _06211_ net65 VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__a21oi_1
X_13585_ _04489_ net694 net757 VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__nand3_1
XFILLER_40_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12536_ _03194_ _03197_ _03332_ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__nand3_1
X_19092_ _09166_ _09384_ _09978_ _09980_ VGND VGND VPWR VPWR _09983_ sky130_fd_sc_hd__o22a_1
XFILLER_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18043_ _08853_ _08888_ _08889_ VGND VGND VPWR VPWR _08893_ sky130_fd_sc_hd__nand3b_1
X_12467_ net679 net483 VGND VGND VPWR VPWR _03399_ sky130_fd_sc_hd__nand2_1
X_15255_ net722 net837 a_h\[12\] net726 VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11418_ net658 net539 VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__nand2_1
X_14206_ _05109_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__inv_2
X_15186_ _05996_ _06051_ _06049_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__a21oi_1
XFILLER_141_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_125_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12398_ _03327_ _03328_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__nand3_4
X_14137_ net724 net709 net703 net728 VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_111_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11349_ _02288_ _02289_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__nand2_1
XFILLER_99_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19994_ net742 net553 VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nand2_1
X_18945_ _09831_ _09825_ _09797_ _09833_ VGND VGND VPWR VPWR _09837_ sky130_fd_sc_hd__o211ai_4
X_14068_ net761 net667 VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__nand2_1
X_13019_ _03938_ _03939_ _03941_ _03799_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a22o_1
X_18876_ _09742_ _09762_ _09763_ _09740_ VGND VGND VPWR VPWR _09768_ sky130_fd_sc_hd__a31o_1
X_17827_ net900 net473 VGND VGND VPWR VPWR _08688_ sky130_fd_sc_hd__nand2_1
XFILLER_81_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17758_ _08619_ net137 VGND VGND VPWR VPWR _08621_ sky130_fd_sc_hd__nor2_1
X_16709_ _07578_ _07580_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__nand2_1
XFILLER_81_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17689_ _08550_ _08551_ VGND VGND VPWR VPWR _08552_ sky130_fd_sc_hd__nand2_1
XFILLER_62_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19428_ net603 net725 VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__nand2_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19359_ _00491_ _00533_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__nand2_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold410 p_hh_pipe\[9\] VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap140 _01630_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xhold443 p_hh_pipe\[8\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap151 _02442_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xhold432 p_hh\[7\] VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 p_ll_pipe\[11\] VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap162 _06334_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_1
X_20203_ net181 _01442_ _01444_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold421 p_ll_pipe\[25\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 p_hh_pipe\[16\] VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 p_hh\[19\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap173 _06729_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_6
Xhold465 p_ll_pipe\[30\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap195 _04967_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_129_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold498 term_low\[14\] VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20134_ net1013 net728 net557 net724 VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__nand4_1
XFILLER_98_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20065_ net735 net551 net549 net742 VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__a22oi_4
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10720_ _01752_ _01751_ net796 VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10651_ _01691_ _01692_ _01694_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10582_ net795 net1187 VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__and2_1
XFILLER_127_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13370_ _04220_ _04223_ _04224_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_62_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12321_ _03132_ _03133_ _03129_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__a21oi_1
XFILLER_119_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12252_ _03054_ _03184_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__nand2_1
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15040_ _05933_ _05935_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__o21ai_1
X_11203_ _02055_ _02056_ _01992_ _01993_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__o211ai_2
XFILLER_123_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12183_ _02688_ net147 _02959_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__o21a_1
XFILLER_123_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16991_ _07850_ _07852_ _07860_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__nand3_1
X_11134_ _01962_ _02004_ _02008_ _02003_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__a22oi_2
XFILLER_135_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15942_ _06808_ _06809_ _06784_ _06787_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__o211ai_2
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11065_ _01962_ _02004_ _02007_ _01857_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__o2bb2ai_2
X_18730_ _09144_ _09308_ _04555_ _06521_ VGND VGND VPWR VPWR _09616_ sky130_fd_sc_hd__o22a_1
XFILLER_88_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18661_ _09538_ _09539_ net1128 net732 VGND VGND VPWR VPWR _09541_ sky130_fd_sc_hd__nand4_1
XFILLER_49_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15873_ _06689_ _06704_ _06691_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__a21boi_1
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17612_ _08470_ _08471_ net414 VGND VGND VPWR VPWR _08476_ sky130_fd_sc_hd__and3_1
X_18592_ _09199_ _09210_ net457 _09264_ _09188_ VGND VGND VPWR VPWR _09465_ sky130_fd_sc_hd__o32a_1
X_14824_ _05613_ _05614_ _05617_ _05612_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__a22o_1
X_11967_ _02735_ _02899_ net644 net535 _02898_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__o2111ai_4
X_17543_ _08405_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__nand2_1
XFILLER_44_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14755_ net163 _05652_ _05538_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__nand3_1
X_10918_ net713 net530 VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__and2_1
X_17474_ _08230_ _08235_ _08338_ VGND VGND VPWR VPWR _08340_ sky130_fd_sc_hd__nand3_1
XFILLER_60_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13706_ net456 _04610_ net762 net683 VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__and4b_1
X_16425_ net281 _07166_ _07164_ _07161_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__o2bb2ai_1
X_11898_ net682 net497 net492 net687 VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__a22oi_2
X_19213_ _10104_ _10106_ _10074_ VGND VGND VPWR VPWR _10110_ sky130_fd_sc_hd__a21o_1
X_14686_ _05581_ _05583_ _05566_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__a21o_1
X_10849_ net793 net1261 VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__and2_1
X_13637_ _04536_ _04542_ _04544_ _04503_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__o211ai_4
X_16356_ net572 net528 VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__nand2_1
X_13568_ _04382_ net1068 _04474_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__nand3b_4
XFILLER_9_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19144_ net818 net881 net552 net549 VGND VGND VPWR VPWR _10036_ sky130_fd_sc_hd__nand4_4
X_16287_ _07088_ _07155_ _07156_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__nand3_2
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12519_ _03425_ _03444_ _03446_ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__nor3_2
X_19075_ _09957_ _09961_ _09965_ _09962_ VGND VGND VPWR VPWR _09966_ sky130_fd_sc_hd__o211ai_4
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15307_ _06130_ _06135_ _06199_ _06200_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__a22oi_1
X_18026_ _08873_ _08874_ _09155_ _09188_ VGND VGND VPWR VPWR _08876_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13499_ _04406_ _04408_ _04407_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_10_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15238_ _06087_ _06088_ _06128_ _06047_ _06131_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__o221ai_2
XFILLER_126_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15169_ _06058_ _06060_ _06062_ _05897_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19977_ net821 net1102 _09373_ _09264_ VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__a211o_1
X_18928_ _09155_ _09319_ _09658_ _09816_ _09815_ VGND VGND VPWR VPWR _09820_ sky130_fd_sc_hd__o221a_1
XFILLER_95_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18859_ net603 net1091 VGND VGND VPWR VPWR _09751_ sky130_fd_sc_hd__nand2_1
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20752_ clknet_leaf_49_clk _00392_ VGND VGND VPWR VPWR p_ll\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ clknet_leaf_57_clk _00323_ VGND VGND VPWR VPWR p_hl\[17\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_102_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_28_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20117_ _01352_ _01345_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__nand2_1
XFILLER_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20048_ _01200_ _01255_ _01254_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_37_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12870_ _03761_ _03677_ _03760_ _03765_ VGND VGND VPWR VPWR _03798_ sky130_fd_sc_hd__a31o_1
X_11821_ _02754_ _02719_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14540_ net771 net1135 VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__nand2_1
X_11752_ _02560_ _02687_ _02688_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__nand3_1
XFILLER_81_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_37_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _02497_ _02503_ _02500_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__a21oi_2
XFILLER_81_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10703_ p_hl\[11\] p_lh\[11\] _01738_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__o21a_1
X_14471_ _05325_ _05329_ _05364_ _05365_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o2bb2ai_2
X_16210_ _06847_ _07029_ net422 _07084_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__or4b_1
X_10634_ p_hl\[2\] p_lh\[2\] VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__nand2_1
X_17190_ _07923_ _08055_ net571 net503 _08054_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__o2111ai_4
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13422_ _04332_ _04331_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nand2_4
X_16141_ _07014_ _07016_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__nand2_1
X_13353_ _04264_ _04263_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_46_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ _03232_ _03237_ _03233_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__nand3_2
X_10565_ net794 net1277 VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__and2_1
X_10496_ net793 _01649_ _01651_ _01652_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__and4_1
X_16072_ net797 _06947_ _06948_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__nor3_1
X_13284_ _04193_ _04196_ _04192_ VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__o21ai_1
XFILLER_142_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12235_ _03028_ net293 _03165_ _03166_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__nand4_4
XFILLER_6_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15023_ _05808_ _05809_ _05806_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__a21boi_2
X_19900_ _01113_ _01116_ _01119_ _01115_ VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__o211ai_2
XFILLER_30_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12166_ net177 _03089_ net199 _03088_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__o211a_1
XFILLER_122_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19831_ _00996_ _00998_ _01044_ _01045_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__o211ai_2
X_11117_ _02057_ _02058_ _02059_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__o21a_1
XFILLER_111_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16974_ _07775_ _07776_ _07840_ _07779_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__a22oi_1
X_12097_ net293 _03027_ _02995_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__a21o_1
XFILLER_96_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19762_ _00710_ _00855_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__nor2_1
X_11048_ _01882_ _01938_ _01989_ _01902_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__nor4_2
X_15925_ _06692_ _06697_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__nand2_1
Xinput8 a[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_18713_ net626 net729 _09351_ _09166_ VGND VGND VPWR VPWR _09597_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19693_ _00759_ _00750_ _00758_ _00764_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__a22oi_4
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15856_ _06644_ _06727_ net173 _06731_ VGND VGND VPWR VPWR _06735_ sky130_fd_sc_hd__nand4_2
X_18644_ _09468_ net302 _09512_ _09518_ VGND VGND VPWR VPWR _09522_ sky130_fd_sc_hd__o211a_1
X_14807_ _05672_ _05704_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__nand2_4
X_15787_ _06659_ _06661_ _06657_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__a21o_1
XFILLER_92_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18575_ _09386_ _09350_ _09392_ VGND VGND VPWR VPWR _09446_ sky130_fd_sc_hd__a21oi_4
X_12999_ _03921_ _03923_ _03924_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a21o_1
X_17526_ _08387_ _08389_ _08388_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__a21o_1
X_14738_ _05596_ _05598_ _05635_ _05637_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__o2bb2ai_4
X_17457_ _09242_ _09668_ _08319_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_15_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14669_ net756 net649 VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__nand2_1
XFILLER_33_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16408_ _07256_ _07257_ _07277_ _07278_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__o2bb2ai_1
X_17388_ _08250_ net472 net606 VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__and3_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16339_ _07206_ _07211_ _07207_ VGND VGND VPWR VPWR _07213_ sky130_fd_sc_hd__and3_1
X_19127_ _10014_ _10015_ VGND VGND VPWR VPWR _10017_ sky130_fd_sc_hd__nand2_1
X_19058_ _09947_ _09948_ VGND VGND VPWR VPWR _09949_ sky130_fd_sc_hd__nor2_1
XFILLER_126_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18009_ net627 net769 VGND VGND VPWR VPWR _08859_ sky130_fd_sc_hd__nand2_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20804_ clknet_leaf_4_clk _00444_ VGND VGND VPWR VPWR b_h\[10\] sky130_fd_sc_hd__dfxtp_4
X_20735_ clknet_leaf_32_clk _00375_ VGND VGND VPWR VPWR p_ll\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20666_ clknet_leaf_38_clk _00306_ VGND VGND VPWR VPWR p_hl\[0\] sky130_fd_sc_hd__dfxtp_1
Xwire428 _05477_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20597_ clknet_leaf_14_clk _00237_ VGND VGND VPWR VPWR p_hh_pipe\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10350_ _01106_ _01161_ _01095_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__o21bai_1
X_10281_ term_low\[19\] term_mid\[19\] VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__nand2_1
X_12020_ _02949_ _02952_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__o21ai_1
XFILLER_132_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13971_ net771 net1122 net667 net660 VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__nand4_1
X_16690_ _07486_ _07488_ _07555_ _07557_ VGND VGND VPWR VPWR _07562_ sky130_fd_sc_hd__a22o_1
X_15710_ net595 net1041 net522 net1120 VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__a22oi_2
X_12922_ _03732_ _03839_ _03840_ _03809_ VGND VGND VPWR VPWR _03850_ sky130_fd_sc_hd__a31o_1
XFILLER_58_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15641_ net616 net611 net531 net527 VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__nand4_2
XFILLER_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12853_ _03715_ _03779_ _03780_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__nand3_2
X_15572_ _06450_ _06452_ _06430_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__o21bai_4
X_11804_ _02737_ _02739_ _02733_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a21o_1
X_18360_ _09209_ _09211_ _09212_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__a21boi_1
X_12784_ _03620_ _03622_ _03691_ VGND VGND VPWR VPWR _03713_ sky130_fd_sc_hd__o21ai_1
X_11735_ _02604_ _02670_ _02672_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__nand3_2
X_17311_ net449 _08173_ _08166_ _08172_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__o211ai_2
X_18291_ net769 net604 net1113 net1123 VGND VGND VPWR VPWR _09137_ sky130_fd_sc_hd__a22oi_4
XPHY_EDGE_ROW_54_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14523_ _09264_ _09471_ _05421_ _05422_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__o211ai_2
XFILLER_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17242_ _08104_ _08109_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__nand2_1
XFILLER_42_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14454_ _05336_ _05338_ _05353_ _05354_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_12_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11666_ _02598_ _02601_ _02603_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__o21ai_4
X_13405_ net196 _04313_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__nand2_1
X_11597_ _02532_ _02533_ _02535_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__a21oi_1
X_17173_ _09373_ _09602_ VGND VGND VPWR VPWR _08041_ sky130_fd_sc_hd__nor2_1
X_10617_ net794 net1217 VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__and2_1
X_14385_ net454 _05158_ net1145 _05287_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__o211ai_4
X_10548_ net793 net1265 VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__and2_1
X_16124_ net595 net570 net1063 net521 VGND VGND VPWR VPWR _07000_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_77_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13336_ _04213_ _04214_ _04246_ _04247_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__nand4_1
Xmax_cap706 a_h\[2\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__buf_8
XFILLER_6_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap717 b_l\[15\] VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__buf_8
Xmax_cap728 b_l\[12\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__buf_8
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16055_ _06927_ net238 VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__nand2_4
X_13267_ net953 net710 net704 net923 VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__a22o_1
Xmax_cap739 net740 VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__buf_12
X_10479_ term_mid\[43\] term_high\[43\] _01613_ _01614_ _01639_ VGND VGND VPWR VPWR
+ _01640_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_90_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12218_ net644 net638 net526 net524 VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__nand4_2
X_15006_ _05819_ _05903_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__nand2_1
XFILLER_142_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_63_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13198_ _04096_ _04102_ _04104_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__a21oi_1
X_12149_ _03035_ _03037_ _03081_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__a21oi_4
XFILLER_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19814_ _01025_ _01013_ _01024_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__nand3_2
XFILLER_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16957_ _07818_ _07823_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__nand2_1
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19745_ _00950_ _00949_ _00869_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__nand3_4
X_15908_ _06769_ _06770_ _06776_ _06777_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_65_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16888_ _07753_ _07755_ _09231_ _09646_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_92_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19676_ net880 net819 net556 net552 _00871_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__a41o_1
X_15839_ _06623_ _06630_ _06715_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_88_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18627_ _09220_ _09242_ net805 _06985_ _09501_ VGND VGND VPWR VPWR _09503_ sky130_fd_sc_hd__o221a_1
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18558_ _09323_ _09425_ VGND VGND VPWR VPWR _09429_ sky130_fd_sc_hd__nand2_1
X_17509_ _08228_ _08295_ _08334_ _08335_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__o211ai_4
XANTENNA_13 _00435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18489_ _09232_ _09244_ _09245_ _09259_ _09243_ VGND VGND VPWR VPWR _09353_ sky130_fd_sc_hd__a32oi_4
XFILLER_60_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20520_ clknet_leaf_42_clk _00160_ VGND VGND VPWR VPWR term_low\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_35 net1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20451_ clknet_leaf_17_clk _00091_ VGND VGND VPWR VPWR term_high\[43\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20382_ clknet_leaf_32_clk _00022_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput120 net120 VGND VGND VPWR VPWR p[59] sky130_fd_sc_hd__buf_2
XFILLER_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11520_ net983 net487 _02455_ _02456_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__a22o_1
XFILLER_51_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20718_ clknet_leaf_22_clk _00358_ VGND VGND VPWR VPWR p_lh\[20\] sky130_fd_sc_hd__dfxtp_1
Xwire203 _01265_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__buf_1
Xwire214 _01407_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__buf_1
X_20649_ clknet_leaf_15_clk _00289_ VGND VGND VPWR VPWR p_hh\[15\] sky130_fd_sc_hd__dfxtp_1
X_11451_ _02291_ _02295_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__nand2_1
XFILLER_7_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10402_ term_mid\[37\] term_high\[37\] VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__and2_1
X_11382_ _02240_ _02319_ _02320_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__nand3_2
X_14170_ _05073_ _05074_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_59_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13121_ a_h\[13\] b_h\[14\] _04042_ _04043_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__a22o_1
X_10333_ term_low\[27\] term_mid\[27\] VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__xor2_1
XFILLER_127_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10264_ term_low\[16\] net1316 net797 VGND VGND VPWR VPWR _10029_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_72_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13052_ net1015 net976 net463 _03896_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__a31o_1
X_12003_ _02788_ _02791_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__nand2_1
X_17860_ _08719_ net477 net1006 _08718_ VGND VGND VPWR VPWR _08720_ sky130_fd_sc_hd__and4_1
X_10195_ b_l\[11\] VGND VGND VPWR VPWR _09308_ sky130_fd_sc_hd__inv_16
XFILLER_120_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16811_ _09242_ _09613_ _07353_ _07498_ VGND VGND VPWR VPWR _07682_ sky130_fd_sc_hd__o22a_1
XFILLER_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17791_ _08554_ _08557_ _08580_ _08583_ _08649_ VGND VGND VPWR VPWR _08653_ sky130_fd_sc_hd__o221ai_4
Xclone126 net924 VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__clkbuf_16
X_19530_ net887 net717 VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__nand2_1
X_16742_ _09210_ _09646_ _02338_ _06761_ _07608_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__o221ai_2
XFILLER_47_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13954_ _04608_ _04720_ _04722_ _04718_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__o22ai_2
X_16673_ _07511_ _07542_ _07543_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__and3_1
X_12905_ _03828_ _03829_ _09504_ _09646_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_46_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13885_ _09177_ _09329_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__nor2_1
X_19461_ _10166_ _10167_ _10171_ _10165_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__a22o_1
X_15624_ net632 net512 VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__nand2_1
X_12836_ _03631_ _03633_ _03652_ _03654_ VGND VGND VPWR VPWR _03765_ sky130_fd_sc_hd__a31o_1
X_18412_ net1100 net749 VGND VGND VPWR VPWR _09269_ sky130_fd_sc_hd__and2_1
X_19392_ _10152_ _00573_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__nand2_1
X_15555_ net625 net532 VGND VGND VPWR VPWR _06438_ sky130_fd_sc_hd__nand2_1
X_18343_ net276 _09192_ VGND VGND VPWR VPWR _09194_ sky130_fd_sc_hd__nor2_1
XFILLER_61_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12767_ _03693_ _03613_ _03692_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__nand3_2
X_14506_ _05407_ _05408_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__nand2_1
X_11718_ _09428_ _09613_ _02653_ _02654_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__o211ai_4
X_12698_ net674 net669 b_h\[12\] net481 VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__nand4_2
X_18274_ _09116_ net759 net804 VGND VGND VPWR VPWR _09120_ sky130_fd_sc_hd__nand3_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15486_ _06355_ _06372_ _06373_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__and3_1
XFILLER_128_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11649_ _02585_ _02586_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__nand2_1
X_17225_ _07920_ net343 _07934_ VGND VGND VPWR VPWR _08093_ sky130_fd_sc_hd__a21boi_2
Xinput11 a[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput22 a[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
X_14437_ _05336_ _05338_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__nor2_1
X_17156_ _07728_ _07730_ _07879_ _07881_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__nand4_1
Xinput33 b[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput44 b[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 b[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
X_14368_ net771 net642 VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__nand2_4
X_16107_ _06866_ _06981_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__nand2_2
Xmax_cap525 net526 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_12
Xmax_cap536 b_h\[2\] VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__buf_12
Xmax_cap503 net504 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_8
X_13319_ _04219_ _04226_ _04227_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__nand3_2
Xmax_cap514 b_h\[6\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17087_ _09242_ _09646_ _02338_ _06985_ _07954_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__o221ai_4
Xmax_cap558 net559 VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkbuf_8
Xmax_cap569 a_l\[11\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__buf_12
X_14299_ net730 net695 VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__nand2_1
X_16038_ _06858_ _06888_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__nand2_2
XFILLER_69_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17989_ net781 net615 net611 net790 VGND VGND VPWR VPWR _08840_ sky130_fd_sc_hd__a22oi_4
XFILLER_93_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19728_ _00907_ _00908_ _00932_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__o21ai_2
XFILLER_37_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19659_ _00729_ _00836_ _00835_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__a21boi_2
XFILLER_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20503_ clknet_leaf_16_clk _00143_ VGND VGND VPWR VPWR term_mid\[47\] sky130_fd_sc_hd__dfxtp_1
XFILLER_119_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20434_ clknet_leaf_15_clk _00074_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfxtp_1
X_20365_ clknet_leaf_49_clk _00005_ VGND VGND VPWR VPWR b_l\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20296_ _01521_ _01526_ _01541_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10951_ _01896_ _01897_ _01883_ _01884_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__a211o_1
XFILLER_44_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13670_ _04574_ _04575_ _04475_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nand3_4
X_12621_ _03397_ _03550_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__nand2_1
X_10882_ net794 net1232 VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12552_ _03480_ _03479_ _03482_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__a21o_1
X_15340_ _06227_ _06231_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_42_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _02141_ _02233_ _02328_ _02332_ _02334_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o32a_1
X_12483_ _03411_ _03412_ _03414_ VGND VGND VPWR VPWR _03415_ sky130_fd_sc_hd__a21o_2
X_15271_ _06095_ _06164_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__nand2_1
XFILLER_8_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _07722_ net144 _07718_ _07876_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__o211ai_1
X_11434_ net672 net525 VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__nand2_1
XFILLER_8_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14222_ net750 net667 VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__nand2_1
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11365_ _02288_ _02289_ _02301_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__a21o_1
X_14153_ net740 net917 net695 net690 VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nand4_1
X_11296_ _02237_ _02148_ net796 VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a21oi_1
X_13104_ _03989_ _03957_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__nand2_1
X_18961_ _09851_ _09849_ _09848_ VGND VGND VPWR VPWR _09853_ sky130_fd_sc_hd__nand3b_4
X_14084_ net788 net783 net643 net639 VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__nand4_4
X_10316_ _00795_ _00838_ _00827_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__and3_1
XFILLER_112_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_112_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10247_ net794 net1166 VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__and2_1
X_17912_ _08711_ _08746_ VGND VGND VPWR VPWR _08771_ sky130_fd_sc_hd__nor2_1
X_13035_ _03891_ _03959_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__nand2_1
XFILLER_3_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18892_ net1111 net747 _09779_ _09780_ VGND VGND VPWR VPWR _09784_ sky130_fd_sc_hd__a22o_1
X_17843_ _08701_ _08702_ _08703_ VGND VGND VPWR VPWR _08704_ sky130_fd_sc_hd__a21o_1
X_17774_ a_l\[15\] net494 net490 net555 VGND VGND VPWR VPWR _08636_ sky130_fd_sc_hd__a22o_1
XFILLER_66_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14986_ _05658_ _05775_ _05776_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__a21o_1
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16725_ net843 net477 VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__nand2_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19513_ _09144_ _09384_ _00546_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13937_ net735 net699 net695 net742 VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_85_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19444_ _00624_ _00625_ net297 VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16656_ net533 net558 net566 net529 VGND VGND VPWR VPWR _07528_ sky130_fd_sc_hd__nand4_4
XFILLER_90_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13868_ _04770_ _04765_ _04653_ _04771_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__o211a_1
X_16587_ _07456_ _07457_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__nand2_1
X_15607_ _06474_ _06483_ _06484_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__nand3_1
X_12819_ _03745_ _03746_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__nand2_1
X_19375_ _00551_ _00553_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__nand2_2
X_13799_ net746 net694 VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__nand2_1
X_15538_ _06404_ _06418_ _06420_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__nand3_1
X_18326_ _09126_ _09127_ _09171_ VGND VGND VPWR VPWR _09175_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18257_ net219 _09018_ net188 _09099_ _09097_ VGND VGND VPWR VPWR _09104_ sky130_fd_sc_hd__o2111ai_2
X_15469_ net716 net650 _06321_ _06319_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__a31o_1
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17208_ _08049_ _07907_ _08048_ _08075_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__o211a_1
X_18188_ _08983_ _08986_ _08987_ VGND VGND VPWR VPWR _09035_ sky130_fd_sc_hd__a21oi_2
X_17139_ _08004_ _08005_ net159 VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__a21oi_1
Xmax_cap344 _07656_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_2
Xmax_cap377 _07743_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_2
Xmax_cap355 _03404_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__buf_1
X_20150_ _01388_ net574 _01387_ b_l\[15\] VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__nand4_2
XFILLER_131_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap399 _02831_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_2
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20081_ _01312_ _01313_ _01101_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__a21o_1
Xmax_cap388 _06314_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_1
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_127_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20417_ clknet_leaf_18_clk _00057_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfxtp_1
X_11150_ _02086_ _02090_ _02092_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__o21ai_1
XFILLER_107_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20348_ net794 net45 VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__and2_1
XFILLER_134_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ _02022_ _02023_ _02018_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__and3_1
X_20279_ _01522_ _01523_ _01499_ net141 VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__a22oi_1
XFILLER_75_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14840_ _05621_ _05626_ _05728_ _05734_ _05733_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__o221a_4
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14771_ _05583_ _05565_ _05561_ _05586_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__o211ai_2
X_16510_ _07372_ _07378_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__nand2_1
X_11983_ _02910_ _02915_ _02917_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__o21ai_1
XFILLER_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13722_ _04506_ _04508_ _04509_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__a21oi_2
X_10934_ _01865_ _01880_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__nand2_1
X_17490_ _08348_ _08349_ _08354_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10865_ net793 net1299 VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__and2_1
X_16441_ net841 net484 net480 net629 VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__a22o_1
XFILLER_71_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13653_ _04558_ _04560_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__nor2_1
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16372_ net586 net515 VGND VGND VPWR VPWR _07246_ sky130_fd_sc_hd__nand2_1
X_12604_ net354 _03443_ _03440_ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a21boi_4
XTAP_TAPCELL_ROW_80_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ _04490_ net701 net751 VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__nand3_1
X_19160_ _10049_ _10052_ VGND VGND VPWR VPWR _10053_ sky130_fd_sc_hd__nand2_1
XFILLER_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10796_ _01808_ _01814_ _01806_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__o21bai_1
X_12535_ net696 _03303_ net475 _03301_ VGND VGND VPWR VPWR _03467_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_80_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18111_ _08904_ _08907_ _08909_ _08957_ VGND VGND VPWR VPWR _08959_ sky130_fd_sc_hd__o211a_1
X_15323_ _06216_ _06217_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__nand2_1
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19091_ _09166_ _09384_ VGND VGND VPWR VPWR _09982_ sky130_fd_sc_hd__nor2_1
XFILLER_138_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18042_ _08856_ _08890_ VGND VGND VPWR VPWR _08892_ sky130_fd_sc_hd__nor2_1
X_12466_ net682 net481 VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__nand2_1
X_15254_ net722 net837 net870 net726 VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__a22oi_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12397_ _03138_ _03140_ _03139_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__a21boi_2
X_11417_ net664 net536 VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__nand2_1
X_14205_ _05073_ _05080_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__a21o_1
X_15185_ _06080_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__inv_2
XFILLER_141_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11348_ _02280_ _02281_ _02286_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__nand3_4
X_14136_ _04932_ _04935_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_111_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19993_ net735 net557 VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__nand2_1
XFILLER_140_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11279_ _02115_ _02117_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__and2_1
X_18944_ _09797_ _09833_ VGND VGND VPWR VPWR _09836_ sky130_fd_sc_hd__nand2_1
X_14067_ _04906_ _04970_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__nand2_1
X_13018_ _03942_ _03940_ VGND VGND VPWR VPWR _03945_ sky130_fd_sc_hd__or2_1
X_18875_ _09742_ _09762_ _09763_ VGND VGND VPWR VPWR _09767_ sky130_fd_sc_hd__nand3_2
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17826_ _08672_ _08686_ VGND VGND VPWR VPWR _08687_ sky130_fd_sc_hd__xnor2_1
XFILLER_67_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17757_ _08271_ _08368_ _08615_ VGND VGND VPWR VPWR _08620_ sky130_fd_sc_hd__nor3_2
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14969_ _05864_ _05792_ _05863_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__nand3_4
X_16708_ _07575_ _07576_ _07433_ VGND VGND VPWR VPWR _07580_ sky130_fd_sc_hd__a21o_1
X_17688_ net565 net485 VGND VGND VPWR VPWR _08551_ sky130_fd_sc_hd__nand2_1
X_16639_ net307 _07399_ _07389_ VGND VGND VPWR VPWR _07511_ sky130_fd_sc_hd__a21boi_1
X_19427_ net887 net718 VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__nand2_1
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19358_ _00488_ _00490_ _00532_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__a21oi_2
X_18309_ _09155_ _09242_ _09150_ _09151_ VGND VGND VPWR VPWR _09157_ sky130_fd_sc_hd__o211ai_1
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19289_ net1148 net579 _00458_ _00460_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__a22o_4
Xhold400 term_low\[13\] VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 p_ll\[18\] VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 p_hh_pipe\[2\] VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap130 _08670_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xhold433 p_ll_pipe\[12\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 p_ll\[17\] VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
X_20202_ _01438_ net182 net214 VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__o21bai_1
XFILLER_145_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold466 p_hh\[14\] VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 mid_sum\[16\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap196 net197 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
Xhold455 p_ll_pipe\[14\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 p_hh\[6\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 p_hh\[27\] VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20133_ net563 net728 net557 VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__nand3_1
XFILLER_58_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_51_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20064_ net742 net549 VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ p_hl\[3\] p_lh\[3\] _01690_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__a21oi_1
XFILLER_41_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10581_ net795 net1195 VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_108_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12320_ _09471_ _09613_ _03129_ _03131_ _02976_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__o32a_2
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12251_ net1048 net995 net492 net679 VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__a22oi_1
X_11202_ _02060_ net180 _02142_ _02143_ _02139_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__a311o_1
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12182_ _02813_ _02962_ _02959_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__o21ai_4
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16990_ _07858_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__nand2_1
X_11133_ _01962_ _02004_ _02008_ _02003_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__a22o_1
X_15941_ _06784_ _06787_ _06813_ _06814_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11064_ net681 net678 net965 net538 VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__nand4_1
X_18660_ net1128 net732 _09538_ _09539_ VGND VGND VPWR VPWR _09540_ sky130_fd_sc_hd__a22o_1
X_15872_ _06704_ _06689_ _06684_ _06690_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__o2bb2ai_2
X_17611_ _08470_ _08471_ net414 VGND VGND VPWR VPWR _08475_ sky130_fd_sc_hd__a21o_1
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18591_ _09450_ _09457_ _09458_ VGND VGND VPWR VPWR _09464_ sky130_fd_sc_hd__nand3_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14823_ _05718_ _05719_ net730 net670 VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__nand4_2
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11966_ _02898_ _02900_ _09515_ _09592_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__o2bb2ai_2
X_17542_ _08404_ _08392_ _08403_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__nand3_1
X_14754_ _05652_ _05538_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__nand2_1
X_10917_ net796 _01864_ _01865_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__nor3_1
X_17473_ _08337_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__nand2_1
XFILLER_44_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13705_ net924 net768 net675 net673 _04607_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__a41o_1
X_14685_ _05580_ _05584_ _05582_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__o21ai_2
X_16424_ _07289_ _07292_ _07294_ VGND VGND VPWR VPWR _07298_ sky130_fd_sc_hd__nand3_1
X_11897_ net682 net499 VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__nand2_1
X_13636_ _04543_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__nand2_1
X_19212_ _10104_ _10106_ _10074_ VGND VGND VPWR VPWR _10109_ sky130_fd_sc_hd__a21oi_1
X_10848_ net793 net1242 VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__and2_1
X_16355_ net561 net541 VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__nand2_1
X_10779_ _01792_ _01799_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__or3_1
X_13567_ _04382_ _04476_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__nand2_2
XFILLER_13_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19143_ net1067 b_l\[2\] net552 net549 VGND VGND VPWR VPWR _10035_ sky130_fd_sc_hd__and4_1
XFILLER_145_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16286_ _07088_ _07155_ _07156_ VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__and3_1
XFILLER_118_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12518_ _03421_ _03423_ _03444_ _03446_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__o22ai_1
X_13498_ net763 net694 _04404_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and3_1
X_19074_ _09794_ _09835_ _09836_ _09832_ VGND VGND VPWR VPWR _09965_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15306_ _06130_ _06135_ _06199_ _06200_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__nand4_2
X_12449_ _03295_ _03378_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__nand2_1
X_18025_ _08873_ _08874_ net779 net615 VGND VGND VPWR VPWR _08875_ sky130_fd_sc_hd__nand4_4
X_15237_ _06132_ _06089_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__nand2_1
XFILLER_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15168_ _05897_ _06062_ _06060_ _06058_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__o211ai_1
X_19976_ _00872_ net548 net895 VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__and3_1
X_14119_ _05021_ _05022_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__nand2_1
X_15099_ _05994_ _05995_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__and2_1
X_18927_ _09817_ net1084 net780 VGND VGND VPWR VPWR _09819_ sky130_fd_sc_hd__nand3_2
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18858_ net609 net737 VGND VGND VPWR VPWR _09750_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_124_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17809_ _08670_ _08669_ net796 VGND VGND VPWR VPWR _08671_ sky130_fd_sc_hd__a21oi_1
XFILLER_55_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18789_ net597 net1001 VGND VGND VPWR VPWR _09681_ sky130_fd_sc_hd__nand2_1
XFILLER_36_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20751_ clknet_leaf_47_clk _00391_ VGND VGND VPWR VPWR p_ll\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_36_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20682_ clknet_leaf_57_clk _00322_ VGND VGND VPWR VPWR p_hl\[16\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_102_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20116_ _01350_ _01351_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__nand2_1
X_20047_ _01189_ _01260_ _01261_ _01265_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__a31o_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11820_ _02717_ _02718_ _02752_ _02753_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__nand4_2
X_11751_ _02687_ _02688_ _02560_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10702_ _01724_ _01728_ _01732_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__nand3_1
XFILLER_53_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _02497_ _02503_ _02500_ VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__a21o_1
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14470_ _05366_ _05370_ _05180_ _05324_ _05329_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__o221ai_4
X_10633_ _01678_ _01675_ _09690_ _01679_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__o211a_1
X_13421_ _04326_ _04328_ _04261_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__o21ai_4
XFILLER_10_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16140_ _07010_ _06976_ _07009_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__nand3_2
X_13352_ _04236_ _04234_ _04237_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__a21o_1
X_10564_ net794 net1272 VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__and2_1
X_16071_ _06845_ _06945_ _06946_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__and3_1
XFILLER_127_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12303_ net177 _03089_ _03098_ _03088_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__a2bb2oi_2
X_10495_ _01651_ _01652_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__nand2_2
X_13283_ net787 net784 net693 net986 VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__nand4_1
X_15022_ _05844_ _05833_ _05834_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__a21boi_2
X_12234_ _03142_ _03143_ _03162_ _03163_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__nand4_1
X_12165_ _03096_ _03097_ _03084_ _03089_ _03088_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_75_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19830_ _01036_ _01037_ _01038_ _00930_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__o2bb2ai_1
X_11116_ _02055_ _02056_ _01991_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__o21ai_2
XFILLER_122_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19761_ _00708_ _00852_ _00854_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__o21ai_1
XFILLER_110_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16973_ _07779_ _07838_ _07839_ VGND VGND VPWR VPWR _07843_ sky130_fd_sc_hd__nand3_4
X_12096_ net293 _03027_ _02995_ VGND VGND VPWR VPWR _03031_ sky130_fd_sc_hd__a21oi_2
X_18712_ net1128 net630 _05043_ VGND VGND VPWR VPWR _09596_ sky130_fd_sc_hd__and3_1
X_11047_ _01934_ _01937_ _01987_ _01988_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__nand4_1
X_15924_ _06798_ _06791_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__nand2_1
X_19692_ _00894_ _00895_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__nand2_2
X_15855_ _06642_ _06564_ _06732_ _06730_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__o211ai_2
X_18643_ _09468_ net302 _09518_ VGND VGND VPWR VPWR _09521_ sky130_fd_sc_hd__o21ai_1
Xinput9 a[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18574_ _09350_ _09386_ _09388_ _09391_ VGND VGND VPWR VPWR _09445_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14806_ net312 _05671_ _05702_ _05703_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__nand4_4
X_15786_ _09166_ _09613_ _06659_ _06661_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__o211ai_1
X_17525_ _08387_ _08389_ _08388_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__a21oi_1
X_12998_ _03921_ _03923_ _03924_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__nand3_2
X_11949_ net647 net526 net1059 net653 VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__a22oi_4
XFILLER_60_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14737_ _05632_ _05599_ _05629_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__nand3_2
X_17456_ _09242_ _09668_ _08319_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_15_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net745 net662 VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__nand2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16407_ _07256_ _07257_ _07273_ _07275_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__o2bb2ai_1
X_17387_ _08247_ _08248_ _08252_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__and3_1
X_13619_ _04349_ _04416_ _04420_ _04414_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__o22a_1
X_16338_ net345 _07210_ _07209_ _07208_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__o211ai_4
X_14599_ _05494_ _05495_ _05496_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__nand3_1
X_19126_ net755 net579 net575 net760 VGND VGND VPWR VPWR _10016_ sky130_fd_sc_hd__a22oi_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_779 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16269_ _07142_ net345 _07138_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__nor3_1
XFILLER_133_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19057_ _09941_ _09943_ _09939_ VGND VGND VPWR VPWR _09948_ sky130_fd_sc_hd__a21oi_2
XFILLER_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18008_ net630 net764 VGND VGND VPWR VPWR _08858_ sky130_fd_sc_hd__nand2_1
XFILLER_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19959_ _00968_ _00969_ _01079_ _01080_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__nand4_2
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20803_ clknet_leaf_4_clk _00443_ VGND VGND VPWR VPWR b_h\[9\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_104_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ clknet_leaf_33_clk _00374_ VGND VGND VPWR VPWR p_ll\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_24_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20665_ clknet_leaf_1_clk _00305_ VGND VGND VPWR VPWR p_hh\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire407 _00733_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_2
Xwire429 _05157_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_2
X_20596_ clknet_leaf_14_clk _00236_ VGND VGND VPWR VPWR p_hh_pipe\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10280_ term_low\[19\] term_mid\[19\] VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__or2_1
XFILLER_132_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone308 net545 VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__clkbuf_16
X_13970_ net771 net767 net667 net660 VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__and4_2
X_12921_ _03732_ _03839_ _03840_ _03809_ VGND VGND VPWR VPWR _03849_ sky130_fd_sc_hd__a31oi_4
XFILLER_58_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15640_ net616 net612 VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__nand2_8
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12852_ _03715_ _03779_ _03780_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__and3_1
XFILLER_33_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15571_ _06430_ _06451_ _06453_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__nand3_1
X_11803_ _02733_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__nand2_2
X_12783_ _03711_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_53_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_8
X_11734_ _02646_ _02666_ net227 _02665_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__o211ai_4
X_17310_ _08174_ net449 _08167_ _08175_ VGND VGND VPWR VPWR _08177_ sky130_fd_sc_hd__o211ai_4
X_18290_ net774 net769 net604 net599 VGND VGND VPWR VPWR _09136_ sky130_fd_sc_hd__nand4_1
XPHY_EDGE_ROW_1_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14522_ _09482_ _09493_ _04260_ _05418_ _05421_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_32_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _02599_ _02600_ net326 VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a21o_1
X_17241_ net582 net573 net498 net493 VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__nand4_2
X_14453_ _05355_ _05340_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13404_ _04174_ _04209_ _04253_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__nor3b_1
X_10616_ net794 net1213 VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__and2_1
XFILLER_128_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11596_ _02393_ _02396_ _02398_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__a21oi_1
X_17172_ _08037_ _08039_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_77_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14384_ _04988_ _05285_ _05284_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__o21ai_1
X_10547_ net793 net1264 VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__and2_1
X_16123_ net570 net522 VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__nand2_2
Xmax_cap707 net708 VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_77_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _04213_ _04214_ _04246_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__a22o_1
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10478_ term_mid\[47\] term_high\[47\] _01637_ _01638_ VGND VGND VPWR VPWR _01639_
+ sky130_fd_sc_hd__a211o_1
X_16054_ _06853_ _06926_ _06927_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__nand3b_4
X_13266_ _04159_ _04169_ _04168_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__o21a_1
Xrebuffer190 _09851_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd1_1
Xmax_cap729 b_l\[12\] VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_90_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12217_ net637 net524 VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__nand2_4
X_15005_ _05820_ _05857_ _05858_ VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__nand3_2
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13197_ net641 net634 b_h\[14\] b_h\[15\] _04117_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__a41o_1
X_19813_ _09286_ _09308_ _00915_ _01020_ _01019_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__o221ai_1
X_12148_ _03035_ _03037_ _03073_ _03075_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__o2bb2ai_4
X_16956_ _07652_ _07816_ _07823_ _07815_ VGND VGND VPWR VPWR _07826_ sky130_fd_sc_hd__o211ai_2
XFILLER_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12079_ _03011_ net518 net906 _03009_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__and4_1
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19744_ _00896_ _00944_ _00945_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__nand3_1
X_15907_ _06778_ _06780_ _06769_ _06770_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__o211ai_2
X_19675_ _00875_ _00877_ _09264_ _09319_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16887_ _07753_ _07755_ _07749_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__a21o_1
XFILLER_65_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18626_ net775 net1131 net589 net581 VGND VGND VPWR VPWR _09502_ sky130_fd_sc_hd__nand4_2
X_15838_ _06711_ _06672_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_88_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15769_ _06504_ _06568_ _06570_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__nand3b_1
X_18557_ _09402_ _09403_ _09422_ VGND VGND VPWR VPWR _09427_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_44_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_8
X_17508_ _08342_ _08346_ _08347_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__a21bo_2
X_18488_ _09233_ _09240_ _09241_ _09254_ _09256_ VGND VGND VPWR VPWR _09352_ sky130_fd_sc_hd__a32oi_4
XFILLER_21_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_14 _00435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ net569 net493 VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__nand2_1
XANTENNA_25 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_20450_ clknet_leaf_17_clk _00090_ VGND VGND VPWR VPWR term_high\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20381_ clknet_leaf_32_clk _00021_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfxtp_1
X_19109_ _09998_ _09999_ VGND VGND VPWR VPWR _10000_ sky130_fd_sc_hd__nand2b_1
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput110 net110 VGND VGND VPWR VPWR p[4] sky130_fd_sc_hd__buf_2
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput121 net121 VGND VGND VPWR VPWR p[5] sky130_fd_sc_hd__buf_2
XFILLER_99_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_8
X_20717_ clknet_leaf_20_clk _00357_ VGND VGND VPWR VPWR p_lh\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20648_ clknet_leaf_15_clk _00288_ VGND VGND VPWR VPWR p_hh\[14\] sky130_fd_sc_hd__dfxtp_1
Xwire237 _07424_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_1
XFILLER_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire248 _02755_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_2
X_11450_ _02385_ _02386_ _02387_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__nand3_2
Xwire215 _01390_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__buf_1
X_10401_ term_mid\[37\] term_high\[37\] VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nor2_1
X_20579_ clknet_leaf_17_clk _00219_ VGND VGND VPWR VPWR p_hh_pipe\[9\] sky130_fd_sc_hd__dfxtp_1
X_11381_ _02241_ _02317_ _02318_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_59_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13120_ _04043_ b_h\[14\] net908 _04042_ VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__nand4_1
X_10332_ net794 _01010_ _01021_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__and3_1
X_13051_ _09482_ _09679_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__nor2_1
X_12002_ net712 net475 _02763_ _02764_ VGND VGND VPWR VPWR _02938_ sky130_fd_sc_hd__a31o_1
XFILLER_105_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10263_ term_low\[16\] term_mid\[16\] VGND VGND VPWR VPWR _10018_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_72_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10194_ net901 VGND VGND VPWR VPWR _09297_ sky130_fd_sc_hd__inv_8
XFILLER_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16810_ _07666_ _07673_ _07675_ VGND VGND VPWR VPWR _07681_ sky130_fd_sc_hd__nand3_2
X_17790_ _08586_ _08650_ _08648_ VGND VGND VPWR VPWR _08652_ sky130_fd_sc_hd__nand3_1
X_16741_ _07609_ _07602_ VGND VGND VPWR VPWR _07612_ sky130_fd_sc_hd__nand2_1
Xclone127 net775 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__clkbuf_16
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13953_ _04855_ _04838_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__nand2_1
X_16672_ _07519_ _07539_ _07510_ VGND VGND VPWR VPWR _07544_ sky130_fd_sc_hd__a21oi_1
X_12904_ _09504_ _09646_ _03826_ _09635_ _03829_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__o221ai_2
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19460_ _10166_ _10167_ _10171_ _10165_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__a22oi_2
X_13884_ _04787_ _04789_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__nand3b_2
X_15623_ _06426_ _06456_ _06502_ _06503_ _09690_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__o311a_1
X_18411_ _09134_ _09137_ _09136_ VGND VGND VPWR VPWR _09268_ sky130_fd_sc_hd__o21ai_1
X_12835_ _03631_ _03633_ _03652_ VGND VGND VPWR VPWR _03764_ sky130_fd_sc_hd__and3_1
XFILLER_61_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19391_ _10005_ _10153_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__nand2_1
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
X_15554_ net1120 net540 VGND VGND VPWR VPWR _06437_ sky130_fd_sc_hd__and2_1
X_18342_ _09187_ _09189_ VGND VGND VPWR VPWR _09193_ sky130_fd_sc_hd__nand2_1
X_12766_ _03577_ _03590_ _03694_ _03695_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__o211ai_4
X_14505_ _05403_ _05264_ _05402_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__nand3b_4
XFILLER_147_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11717_ _02652_ net501 net687 _02651_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__nand4_4
X_12697_ net674 net944 b_h\[12\] net481 VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__and4_1
X_18273_ _09116_ _09117_ VGND VGND VPWR VPWR _09119_ sky130_fd_sc_hd__nand2_1
X_15485_ _06374_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__inv_2
X_11648_ _02581_ net1021 _02577_ _02582_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__o211ai_4
Xinput12 a[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_17224_ _07920_ _07935_ _07933_ _07928_ VGND VGND VPWR VPWR _08092_ sky130_fd_sc_hd__o2bb2ai_2
X_14436_ b_l\[14\] net703 _05332_ _05334_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__a22o_1
X_17155_ _07726_ _07729_ _07879_ _07881_ _07728_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__o2111a_1
Xinput23 a[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
X_11579_ _02487_ _02488_ net359 _02512_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__a22o_1
Xinput45 b[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 b[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_14367_ net761 net655 VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__nand2_2
XFILLER_143_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16106_ net583 net533 net529 net1116 VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__a22oi_4
Xmax_cap504 b_h\[8\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__buf_8
X_13318_ _04229_ _04218_ _04228_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__nand3_1
Xinput56 b[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
XFILLER_115_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap537 net539 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__buf_8
X_17086_ net586 net582 net498 net493 VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__nand4_2
X_14298_ _05055_ _05201_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__nand2_1
Xmax_cap548 net549 VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__buf_8
X_16037_ _06913_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13249_ net787 net784 net700 net693 VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__nand4_1
X_17988_ net790 net781 net615 net611 VGND VGND VPWR VPWR _08839_ sky130_fd_sc_hd__nand4_1
XFILLER_84_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19727_ _00909_ _00910_ _00932_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__o21ai_1
X_16939_ net550 b_h\[2\] VGND VGND VPWR VPWR _07809_ sky130_fd_sc_hd__nand2_1
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19658_ _00729_ _00836_ _00834_ _00829_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18609_ net791 net782 net569 net565 VGND VGND VPWR VPWR _09484_ sky130_fd_sc_hd__nand4_1
XFILLER_53_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19589_ net591 net729 VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_17_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20502_ clknet_leaf_16_clk _00142_ VGND VGND VPWR VPWR term_mid\[46\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20433_ clknet_leaf_15_clk net134 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20364_ clknet_leaf_50_clk _00004_ VGND VGND VPWR VPWR b_l\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_106_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20295_ _01539_ net158 _01525_ _01502_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__o22ai_1
XFILLER_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10950_ _01892_ _01893_ _01894_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_3_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ net794 net1178 VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__and2_1
XFILLER_71_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12620_ net680 net674 net483 net481 VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__nand4_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12551_ _03479_ _03480_ _03482_ VGND VGND VPWR VPWR _03483_ sky130_fd_sc_hd__a21oi_2
X_11502_ net201 _02328_ _02438_ _02441_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o31ai_1
X_12482_ net356 _03322_ _03321_ VGND VGND VPWR VPWR _03414_ sky130_fd_sc_hd__o21a_1
X_15270_ net733 net912 net635 net739 VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__a22oi_2
XFILLER_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ net681 net517 VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_91_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14221_ _05123_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__nand2_2
XFILLER_138_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14152_ net740 net916 net695 net690 VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__and4_1
XFILLER_4_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11364_ _02288_ _02289_ net360 VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__a21oi_1
X_11295_ _02144_ _02236_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__xor2_1
X_13103_ _03981_ _03985_ _04024_ _04025_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__nand4_1
X_18960_ _09846_ _09847_ _09851_ VGND VGND VPWR VPWR _09852_ sky130_fd_sc_hd__nand3_4
X_14083_ net783 net639 VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__nand2_2
X_10315_ _00795_ _00838_ _00827_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__a21o_1
X_17911_ _08766_ _08768_ VGND VGND VPWR VPWR _08770_ sky130_fd_sc_hd__xnor2_2
X_13034_ net976 net645 net1149 net999 VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__nand4_2
X_18891_ _09779_ _09780_ net1111 net747 VGND VGND VPWR VPWR _09783_ sky130_fd_sc_hd__nand4_1
X_10246_ net794 net39 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__and2_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17842_ _09286_ _09679_ _08651_ _08653_ VGND VGND VPWR VPWR _08703_ sky130_fd_sc_hd__o31a_1
XFILLER_67_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17773_ a_l\[15\] net490 VGND VGND VPWR VPWR _08635_ sky130_fd_sc_hd__nand2_1
X_14985_ _05881_ _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__nand2_1
X_16724_ net620 net813 net484 net480 VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__nand4_1
X_19512_ _09144_ _09384_ _00546_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__o21a_1
X_13936_ net740 net695 VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__nand2_2
X_16655_ _07377_ _07525_ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_85_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19443_ net297 _00624_ _00625_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__nand3_4
X_15606_ _06474_ _06484_ VGND VGND VPWR VPWR _06488_ sky130_fd_sc_hd__nand2_1
XFILLER_90_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13867_ _04772_ _04652_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__nand3_4
XFILLER_35_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16586_ a_l\[6\] net496 net491 a_l\[5\] VGND VGND VPWR VPWR _07458_ sky130_fd_sc_hd__a22oi_1
X_12818_ net645 b_h\[9\] b_h\[10\] net648 VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__a22oi_1
X_19374_ _00550_ _00552_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__nor2_1
X_13798_ _04607_ _04610_ _04608_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__a21oi_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15537_ _06417_ _06419_ _06404_ VGND VGND VPWR VPWR _06421_ sky130_fd_sc_hd__o21bai_2
X_12749_ _03676_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__nand2_1
X_18325_ _09131_ _09170_ _09171_ VGND VGND VPWR VPWR _09174_ sky130_fd_sc_hd__nand3_1
X_18256_ _09097_ net189 _09021_ _09099_ VGND VGND VPWR VPWR _09103_ sky130_fd_sc_hd__and4_1
X_15468_ _06324_ net221 _06357_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__nor3_1
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17207_ _08060_ _08065_ _08070_ _08063_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__o211ai_2
X_14419_ _05316_ _05317_ _05297_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__o21ai_2
XFILLER_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18187_ _08984_ _08985_ _08983_ VGND VGND VPWR VPWR _09034_ sky130_fd_sc_hd__o21a_1
Xmax_cap301 _09494_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_4
X_15399_ _06251_ _06290_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__nand2_1
X_17138_ _07850_ _07860_ _07851_ VGND VGND VPWR VPWR _08007_ sky130_fd_sc_hd__a21oi_1
Xmax_cap323 _02906_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__buf_6
Xmax_cap345 _07139_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_96_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap356 _03306_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_1
X_17069_ _07785_ _07919_ _07934_ net343 VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_6_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap389 _05606_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_2
X_20080_ _00872_ _01100_ _01310_ VGND VGND VPWR VPWR _01314_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_139_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_127_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20416_ clknet_leaf_17_clk _00056_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20347_ net794 net43 VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__and2_1
X_11080_ _02022_ _02023_ _02018_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__a21oi_1
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20278_ _01522_ _01523_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__and2_1
XFILLER_103_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14770_ _05598_ _05668_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__nand2_2
X_11982_ _02917_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__inv_2
XFILLER_91_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13721_ _04506_ _04508_ _04509_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__a21o_1
XFILLER_44_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10933_ net713 net707 net441 net364 _01880_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_67_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10864_ net793 net1212 VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__and2_1
X_16440_ net625 net484 net480 net628 VGND VGND VPWR VPWR _07313_ sky130_fd_sc_hd__a22oi_1
XFILLER_71_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13652_ _04556_ _04557_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__o21a_1
X_16371_ net583 net559 net544 net523 VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__nand4_2
X_10795_ _01816_ _01817_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__nor2_1
X_12603_ _03532_ _03533_ VGND VGND VPWR VPWR _03534_ sky130_fd_sc_hd__nand2_1
X_13583_ _01888_ _04260_ net748 net705 _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__o2111ai_4
X_12534_ net696 net474 VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18110_ _08904_ _08907_ _08909_ VGND VGND VPWR VPWR _08958_ sky130_fd_sc_hd__o21a_1
X_19090_ _05044_ _06441_ net411 _09766_ _09768_ VGND VGND VPWR VPWR _09981_ sky130_fd_sc_hd__o2111ai_2
X_15322_ _06214_ _05889_ _05888_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__nand3_4
X_18041_ _08853_ _08856_ _08890_ VGND VGND VPWR VPWR _08891_ sky130_fd_sc_hd__nand3_1
XFILLER_8_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12465_ net680 net481 VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__nand2_1
X_15253_ _06147_ _06148_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__nor2_1
XFILLER_125_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11416_ net664 net536 VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__and2_1
X_12396_ _03126_ _03136_ _03137_ _03139_ _03141_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__a32oi_4
X_15184_ net715 _05993_ net680 _05991_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__a31o_1
X_14204_ _09329_ _09351_ _01860_ _05042_ _05047_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__o32a_1
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11347_ _02282_ _02284_ _02287_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__nand3_2
X_19992_ net742 net735 net557 net1102 VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__nand4_1
X_14135_ _04921_ _04928_ _04929_ _04933_ _04918_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__a32oi_4
XFILLER_141_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11278_ net712 net975 VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__nand2_1
X_18943_ _09796_ _09829_ _09830_ VGND VGND VPWR VPWR _09835_ sky130_fd_sc_hd__nand3_2
X_14066_ _04887_ _04905_ _04904_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__o21ai_1
XFILLER_121_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10229_ net473 VGND VGND VPWR VPWR _09679_ sky130_fd_sc_hd__clkinv_16
X_13017_ _03938_ _03939_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__and3_1
X_18874_ _09765_ _09741_ _09764_ VGND VGND VPWR VPWR _09766_ sky130_fd_sc_hd__nand3_4
X_17825_ _08684_ _08685_ VGND VGND VPWR VPWR _08686_ sky130_fd_sc_hd__nand2_1
X_17756_ _08615_ _08459_ _08617_ VGND VGND VPWR VPWR _08619_ sky130_fd_sc_hd__o21bai_4
XFILLER_48_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16707_ _07433_ _07575_ _07576_ _07434_ _07441_ VGND VGND VPWR VPWR _07579_ sky130_fd_sc_hd__a32oi_1
X_14968_ _05793_ _05861_ _05862_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__nand3_2
X_17687_ a_l\[11\] net479 VGND VGND VPWR VPWR _08550_ sky130_fd_sc_hd__nand2_1
X_13919_ _04693_ _04822_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__nor2_1
X_14899_ net756 net750 net642 net640 VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__and4_1
XFILLER_35_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16638_ _07399_ _07387_ _07380_ _07388_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_90_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19426_ _00608_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__inv_2
XFILLER_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16569_ net795 _07440_ _07441_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__and3_2
X_19357_ _00488_ _00490_ _00530_ _00531_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__nand4_2
XFILLER_16_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18308_ _09152_ _09153_ VGND VGND VPWR VPWR _09156_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_98_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19288_ net896 net579 VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__nand2_1
XFILLER_31_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18239_ _09084_ net277 VGND VGND VPWR VPWR _09086_ sky130_fd_sc_hd__nand2_1
Xhold401 p_ll\[25\] VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 p_hh\[13\] VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 mid_sum\[25\] VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 p_hh\[8\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap153 _09207_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_4
Xmax_cap142 _04831_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xhold423 p_ll_pipe\[15\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__dlygate4sd3_1
X_20201_ net181 _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__nor2_1
Xhold467 p_hh_pipe\[18\] VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap175 _03858_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
Xhold478 p_ll_pipe\[10\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 p_ll\[14\] VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap164 _04817_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
X_20132_ net728 net557 VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__nand2_2
XFILLER_132_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_129_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold489 mid_sum\[6\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20063_ net742 net734 net551 net549 VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__nand4_4
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_142_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_107_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10580_ net795 net1304 VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_62_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12250_ net1048 net995 VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__nand2_1
X_11201_ _02055_ _02056_ _01991_ _02137_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__o211ai_2
X_12181_ _03114_ _03115_ VGND VGND VPWR VPWR _03116_ sky130_fd_sc_hd__and2_1
XFILLER_134_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11132_ net1062 _02007_ _02003_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15940_ _06784_ net283 _06787_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__nand3_1
X_11063_ net681 net678 VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__nand2_1
XFILLER_89_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15871_ _06709_ _06712_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__nand2_1
XFILLER_88_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17610_ _08470_ _08471_ net414 VGND VGND VPWR VPWR _08474_ sky130_fd_sc_hd__a21oi_1
X_14822_ _05718_ _05719_ _09308_ _09460_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__o2bb2ai_1
X_18590_ _09450_ _09457_ _09458_ VGND VGND VPWR VPWR _09463_ sky130_fd_sc_hd__and3_1
XFILLER_45_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11965_ _02898_ _02900_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__nand2_1
X_17541_ _08404_ _08392_ _08403_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__and3_1
X_14753_ _05511_ _05509_ _05510_ net163 _05652_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__o2111ai_1
X_10916_ net364 net441 net707 net713 VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__and4_1
X_17472_ _08297_ _08298_ _08334_ _08335_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__o211ai_2
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ net762 net683 net456 _04609_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__a211oi_1
X_14684_ _05568_ _05578_ _05579_ _05583_ _05565_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__a32oi_4
X_16423_ _07289_ _07292_ _07294_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__a21o_1
X_11896_ _02771_ _02772_ _02775_ _02770_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__a22oi_2
X_13635_ _04539_ _04504_ _04541_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nand3_4
X_19211_ _10076_ _10102_ _10103_ _10073_ VGND VGND VPWR VPWR _10108_ sky130_fd_sc_hd__a31o_1
XFILLER_17_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10847_ net795 net1229 VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__and2_1
X_19142_ _09929_ _09932_ VGND VGND VPWR VPWR _10034_ sky130_fd_sc_hd__nand2_1
X_16354_ _07095_ _07102_ _07098_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__a21oi_1
X_10778_ _01801_ _01802_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__nor2_1
X_13566_ _04472_ _04474_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__nand2_2
X_16285_ _07089_ _07152_ _07153_ net258 _07086_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__a32oi_4
X_12517_ _03422_ _03424_ net322 _03447_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__a22oi_4
X_13497_ net763 net694 _04404_ _04406_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__a22oi_2
X_19073_ _09793_ _09837_ _09834_ _09828_ VGND VGND VPWR VPWR _09964_ sky130_fd_sc_hd__o2bb2ai_1
X_15305_ _06191_ _06198_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__nand2_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12448_ _03298_ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__nand2_1
X_18024_ net790 net781 net886 net605 VGND VGND VPWR VPWR _08874_ sky130_fd_sc_hd__nand4_4
X_15236_ _06130_ _06131_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12379_ net665 net499 net495 net674 VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_93_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15167_ _06061_ _06063_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__nand2_1
XFILLER_141_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19975_ _01194_ _01198_ _01197_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__o21ai_2
X_14118_ _05009_ net981 _05018_ _05019_ _05007_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a32oi_4
X_15098_ _05992_ _05993_ net715 net680 VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__nand4_1
X_14049_ _04952_ _04953_ _04833_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__a21o_1
X_18926_ _09815_ _09817_ _09155_ _09319_ VGND VGND VPWR VPWR _09818_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_39_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18857_ net619 net732 VGND VGND VPWR VPWR _09749_ sky130_fd_sc_hd__nand2_1
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17808_ _08612_ _08621_ _08624_ _08613_ VGND VGND VPWR VPWR _08670_ sky130_fd_sc_hd__o31ai_2
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18788_ net606 net747 VGND VGND VPWR VPWR _09680_ sky130_fd_sc_hd__nand2_1
X_17739_ _08593_ _08598_ _08599_ VGND VGND VPWR VPWR _08602_ sky130_fd_sc_hd__nand3_1
X_20750_ clknet_leaf_43_clk _00390_ VGND VGND VPWR VPWR p_ll\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19409_ _00467_ _00470_ _00469_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__a21boi_1
X_20681_ clknet_leaf_55_clk _00321_ VGND VGND VPWR VPWR p_hl\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20115_ _01184_ _01346_ _01348_ _01347_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__o211ai_4
X_20046_ _01275_ _01276_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__nor2_1
XFILLER_73_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11750_ net178 _02683_ _02552_ _02556_ _02682_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_64_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _01735_ _01736_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__nor2_1
XFILLER_41_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _01857_ _02613_ net652 net535 _02612_ VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__o2111ai_4
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10632_ _01675_ _01677_ p_hl\[0\] net1363 VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__a2bb2o_1
X_13420_ _01855_ _04260_ _04327_ _04329_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__o211ai_2
XFILLER_22_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13351_ net714 net963 net1126 _04262_ VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__a31o_1
X_10563_ net794 net1259 VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__and2_1
X_16070_ _06945_ _06946_ _06845_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__a21oi_1
X_12302_ _03098_ _03088_ net177 _03089_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__o2bb2ai_1
Xrebuffer350 _05873_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__buf_1
X_10494_ term_high\[49\] term_high\[50\] term_high\[51\] _01635_ VGND VGND VPWR VPWR
+ _01652_ sky130_fd_sc_hd__nand4_1
XFILLER_108_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13282_ _04162_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__nor2_1
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15021_ _05844_ _05833_ _05834_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__a21bo_1
XFILLER_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12233_ _03142_ _03143_ _03162_ _03163_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__a22o_1
X_12164_ _03090_ net199 VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_75_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ _01991_ _02055_ _02056_ _01994_ net793 VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__o41a_1
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16972_ _07665_ _07778_ _07835_ _07836_ VGND VGND VPWR VPWR _07842_ sky130_fd_sc_hd__nand4_2
X_12095_ _02991_ _02994_ net293 _03027_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__o211ai_2
X_19760_ _00968_ _00969_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__nand2_1
X_11046_ _01934_ _01937_ _01987_ _01988_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__and4_4
X_15923_ _06658_ _06797_ _06796_ _06792_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__o211ai_1
X_18711_ _09462_ _09467_ _09463_ VGND VGND VPWR VPWR _09595_ sky130_fd_sc_hd__a21oi_2
XFILLER_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19691_ _00771_ net272 _00893_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__nand3b_4
X_15854_ _06644_ _06731_ _06730_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__a21o_1
X_18642_ _09475_ _09513_ _09516_ _09473_ VGND VGND VPWR VPWR _09520_ sky130_fd_sc_hd__a31oi_2
XFILLER_49_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15785_ _06663_ _06655_ _06662_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__nand3_4
XFILLER_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18573_ _09223_ _09431_ _09430_ VGND VGND VPWR VPWR _09444_ sky130_fd_sc_hd__a21boi_1
X_14805_ _05704_ _05672_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__nor2_1
XFILLER_18_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17524_ net1093 net485 _08385_ _08384_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__a31oi_1
X_12997_ _03819_ _03835_ _03837_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__o21ai_2
XFILLER_45_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14736_ _05629_ _05632_ _05599_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__and3_1
XFILLER_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11948_ net1016 net526 VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__nand2_2
X_11879_ _02562_ _02687_ _02688_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__and3_1
X_17455_ _02589_ _06985_ net596 net476 _08318_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__o2111ai_4
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _05271_ _05446_ _05441_ _05444_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__o22a_1
X_16406_ _07277_ _07278_ _07256_ _07257_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__o211ai_1
X_17386_ _08124_ _08245_ _08246_ _08251_ VGND VGND VPWR VPWR _08253_ sky130_fd_sc_hd__a31o_1
XFILLER_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13618_ _04420_ _04414_ _04417_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__o21ai_1
X_14598_ _05495_ _05496_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__nand2_1
X_16337_ net345 _07141_ _07138_ VGND VGND VPWR VPWR _07211_ sky130_fd_sc_hd__o21bai_1
X_13549_ _04437_ _04456_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nand2_1
X_19125_ net753 net579 VGND VGND VPWR VPWR _10015_ sky130_fd_sc_hd__nand2_1
XFILLER_146_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19056_ _09940_ _09946_ VGND VGND VPWR VPWR _09947_ sky130_fd_sc_hd__nor2_2
XFILLER_145_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16268_ _07138_ net345 _07142_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__o21a_1
X_18007_ _08833_ _08846_ _08844_ _08845_ VGND VGND VPWR VPWR _08857_ sky130_fd_sc_hd__o2bb2ai_1
X_16199_ _07065_ _07072_ _07073_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__nand3b_4
XFILLER_126_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15219_ net347 _06106_ _06113_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__o21bai_4
XFILLER_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19958_ _00969_ _01078_ _01080_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__o21ai_4
X_19889_ _01105_ _01107_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__nand2_1
X_18909_ net775 net770 net575 net568 VGND VGND VPWR VPWR _09801_ sky130_fd_sc_hd__nand4_2
XFILLER_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20802_ clknet_leaf_3_clk _00442_ VGND VGND VPWR VPWR b_h\[8\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_104_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20733_ clknet_leaf_35_clk _00373_ VGND VGND VPWR VPWR p_ll\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ clknet_leaf_1_clk _00304_ VGND VGND VPWR VPWR p_hh\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20595_ clknet_leaf_14_clk _00235_ VGND VGND VPWR VPWR p_hh_pipe\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone309 net1108 VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__clkbuf_16
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12920_ _03844_ _03845_ _03808_ VGND VGND VPWR VPWR _03848_ sky130_fd_sc_hd__a21o_1
X_20029_ _01254_ _01256_ _01200_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__a21o_1
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12851_ _03721_ _03724_ _03774_ _03776_ VGND VGND VPWR VPWR _03780_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11802_ net644 net1036 net546 net537 VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nand4_4
XFILLER_15_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15570_ _06447_ _06449_ _06433_ _06434_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__a211o_1
XFILLER_92_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12782_ _03614_ _03618_ _03619_ VGND VGND VPWR VPWR _03711_ sky130_fd_sc_hd__a21bo_1
X_11733_ _02646_ _02666_ net227 _02665_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__o211a_1
XFILLER_42_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14521_ _05422_ _05421_ _05418_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__a21o_1
X_11664_ _02599_ _02600_ net326 VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__nand3_1
X_17240_ _08105_ _08106_ VGND VGND VPWR VPWR _08108_ sky130_fd_sc_hd__nand2_2
X_14452_ net349 _05354_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17171_ _09199_ _09679_ _08035_ _08036_ VGND VGND VPWR VPWR _08039_ sky130_fd_sc_hd__o211ai_1
X_13403_ _04313_ _04314_ _04255_ _04211_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__o2bb2a_1
X_10615_ net794 net1244 VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__and2_1
XFILLER_128_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16122_ net1041 net570 net521 net950 VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__a22o_4
X_11595_ _02396_ net501 net698 VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__and3_1
X_14383_ net783 net778 net1135 net636 VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nand4_4
X_10546_ net793 net1237 VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__and2_1
XFILLER_128_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap708 net710 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_77_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _04200_ _04216_ _04242_ _04243_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__nand4_2
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10477_ term_mid\[47\] term_high\[47\] term_mid\[46\] term_high\[46\] VGND VGND VPWR
+ VPWR _01638_ sky130_fd_sc_hd__o211a_1
X_16053_ _06928_ _06853_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__nand2_1
Xrebuffer191 a_l\[6\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_108_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer180 _07647_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd1_1
X_13265_ _04159_ _04169_ _04168_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__o21ai_1
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12216_ _03007_ _03149_ VGND VGND VPWR VPWR _03150_ sky130_fd_sc_hd__nand2_2
X_15004_ _05900_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13196_ net634 b_h\[15\] _04097_ _04099_ VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__o2bb2a_1
X_19812_ _01023_ _01015_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__nand2_1
X_12147_ _03035_ _03037_ _03074_ _03076_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__nand4_4
XFILLER_69_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16955_ _07819_ _07822_ _07818_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__o21ai_2
XFILLER_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12078_ net906 net518 _03009_ _03011_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__a22o_1
X_19743_ _00894_ _00895_ _00947_ _00948_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__nand4_1
X_15906_ _06751_ _06782_ _06783_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__nand3_2
X_11029_ _01964_ _01969_ _01972_ _01953_ _01952_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__o2111ai_1
X_16886_ _02338_ _06867_ _07749_ VGND VGND VPWR VPWR _07756_ sky130_fd_sc_hd__o21ai_1
XFILLER_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19674_ _00873_ _00874_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__nand2_1
X_15837_ _06668_ _06669_ _06709_ _06710_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__o211ai_2
XFILLER_77_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18625_ _09358_ _09499_ VGND VGND VPWR VPWR _09501_ sky130_fd_sc_hd__nand2_1
XFILLER_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15768_ _06643_ _06645_ _06646_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
X_18556_ _09402_ _09403_ _09419_ _09420_ VGND VGND VPWR VPWR _09426_ sky130_fd_sc_hd__o2bb2ai_2
X_15699_ net628 net512 net505 net632 VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_111_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17507_ _08359_ _08371_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__nand2_1
X_18487_ _09348_ _09349_ VGND VGND VPWR VPWR _09350_ sky130_fd_sc_hd__nand2_2
X_14719_ _05479_ _05616_ net730 net677 _05615_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__o2111ai_1
X_17438_ net578 net488 VGND VGND VPWR VPWR _08304_ sky130_fd_sc_hd__nand2_1
XFILLER_21_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_15 _00435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _05043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17369_ _08201_ _08202_ net234 _08232_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__nand4_1
XFILLER_9_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20380_ clknet_leaf_32_clk _00020_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_118_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19108_ _09996_ _09997_ _09857_ VGND VGND VPWR VPWR _09999_ sky130_fd_sc_hd__nand3_2
Xoutput100 net100 VGND VGND VPWR VPWR p[40] sky130_fd_sc_hd__buf_2
X_19039_ b_l\[0\] net549 VGND VGND VPWR VPWR _09930_ sky130_fd_sc_hd__nand2_1
Xoutput111 net111 VGND VGND VPWR VPWR p[50] sky130_fd_sc_hd__buf_2
Xoutput122 net122 VGND VGND VPWR VPWR p[60] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_132_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_120_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20716_ clknet_leaf_20_clk _00356_ VGND VGND VPWR VPWR p_lh\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20647_ clknet_leaf_15_clk _00287_ VGND VGND VPWR VPWR p_hh\[13\] sky130_fd_sc_hd__dfxtp_1
Xwire227 _02668_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__buf_6
Xwire216 _10127_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
X_10400_ net795 _01571_ _01572_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__and3_1
X_20578_ clknet_leaf_18_clk _00218_ VGND VGND VPWR VPWR p_hh_pipe\[8\] sky130_fd_sc_hd__dfxtp_1
X_11380_ _02319_ _02320_ _02240_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__a21oi_1
Xwire249 _02048_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_59_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10331_ _00956_ _00967_ _00999_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__or3_1
X_10262_ net794 net1334 VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__and2_1
X_13050_ _03958_ _03974_ VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__xnor2_2
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12001_ _02930_ _02926_ _02824_ _02931_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_72_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10193_ net576 VGND VGND VPWR VPWR _09286_ sky130_fd_sc_hd__inv_8
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16740_ _02338_ _06761_ a_l\[5\] net1032 _07608_ VGND VGND VPWR VPWR _07611_ sky130_fd_sc_hd__o2111ai_1
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13952_ _04850_ _04853_ _04839_ _04849_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__o211ai_1
XFILLER_143_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12903_ _03830_ _03822_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__nand2_1
XFILLER_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16671_ _07539_ _07519_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__nand2_1
X_13883_ _04783_ _04784_ _04779_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__a21o_1
X_15622_ _06500_ _06501_ _06458_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__nand3_1
XFILLER_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18410_ _09144_ _09188_ net457 _09123_ VGND VGND VPWR VPWR _09267_ sky130_fd_sc_hd__o31a_1
X_12834_ _03758_ _03755_ _03678_ _03759_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__o211ai_2
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19390_ _00570_ _00571_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__nand2_1
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15553_ _06412_ _06414_ _06415_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__a21oi_1
X_12765_ _03621_ _03623_ _03690_ _03691_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__a22o_1
X_18341_ net457 _06402_ net336 _09038_ _09187_ VGND VGND VPWR VPWR _09192_ sky130_fd_sc_hd__o311a_1
X_11716_ _02524_ net510 net679 VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_83_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ net622 net800 net759 net754 VGND VGND VPWR VPWR _09118_ sky130_fd_sc_hd__nand4_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14504_ _05401_ _05403_ _05264_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__o21bai_4
X_17223_ _07963_ _08088_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__nand2_1
X_12696_ net669 b_h\[12\] VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__nand2_1
XFILLER_70_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15484_ _06372_ _06373_ net222 VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__a21o_1
XFILLER_128_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11647_ _02583_ net1021 _02576_ _02584_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__o211ai_2
X_14435_ _05332_ _05334_ _05335_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__a21oi_2
Xinput13 a[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17154_ _08017_ _08019_ _08021_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__o21ai_1
X_11578_ _02483_ _02489_ _02490_ _02513_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__o211a_1
Xinput46 b[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 b[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 a[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xwire750 net752 VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__buf_12
X_14366_ _05186_ _05236_ _05189_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__a21oi_1
X_10529_ net795 net1184 VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__and2_1
Xmax_cap505 net506 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_8
Xmax_cap527 net529 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_12
X_16105_ net583 net533 VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__nand2_1
X_17085_ _07754_ _07953_ VGND VGND VPWR VPWR _07954_ sky130_fd_sc_hd__nand2_4
X_13317_ _04226_ _04227_ _04219_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__a21oi_1
Xinput57 b[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16036_ _06911_ _06912_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__nand2_4
XFILLER_109_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap538 net539 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_6
X_14297_ _04842_ _05056_ _05052_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__o21ai_1
XFILLER_130_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13248_ net787 net784 net700 net693 VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__and4_1
X_13179_ net634 b_h\[14\] b_h\[15\] net641 VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__a22o_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17987_ net790 net781 net615 net611 VGND VGND VPWR VPWR _08838_ sky130_fd_sc_hd__and4_1
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19726_ _00907_ _00908_ _00927_ _00931_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__o211ai_2
X_16938_ _07641_ _07642_ _07640_ VGND VGND VPWR VPWR _07808_ sky130_fd_sc_hd__a21o_1
X_16869_ net608 net485 VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__nand2_1
X_19657_ _00720_ _00842_ _00846_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__o21ai_2
XFILLER_53_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18608_ net792 net782 net569 net1084 VGND VGND VPWR VPWR _09483_ sky130_fd_sc_hd__and4_1
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19588_ net598 net725 VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__nand2_1
X_18539_ _09216_ _09404_ VGND VGND VPWR VPWR _09408_ sky130_fd_sc_hd__nand2_1
XFILLER_61_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20501_ clknet_leaf_16_clk _00141_ VGND VGND VPWR VPWR term_mid\[45\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20432_ clknet_leaf_15_clk net1357 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20363_ clknet_leaf_50_clk _00003_ VGND VGND VPWR VPWR b_l\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_122_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20294_ _01539_ net158 VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__or2_1
XFILLER_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ net794 net1179 VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__and2_1
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12550_ _03347_ _03354_ _03346_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a21boi_1
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11501_ net201 _02328_ _02439_ _02438_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__o22ai_4
X_12481_ net356 _03322_ _03321_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_22_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _02366_ _02368_ _02355_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__nand3_1
X_14220_ net756 net667 VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__nand2_1
XFILLER_137_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14151_ net736 net690 VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__nand2_2
XFILLER_138_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ _02288_ _02289_ _02302_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__nand3_1
X_13102_ _03981_ _03985_ _04025_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__nand3_1
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11294_ _02235_ net201 _02234_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__a21oi_4
X_14082_ net783 net1135 VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__and2_1
X_10314_ _00698_ _00762_ _00784_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__nand3_1
X_17910_ _08768_ _08766_ VGND VGND VPWR VPWR _08769_ sky130_fd_sc_hd__nor2_1
X_13033_ a_h\[13\] net1149 VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__nand2_1
X_18890_ _09231_ _09264_ _09779_ _09780_ VGND VGND VPWR VPWR _09782_ sky130_fd_sc_hd__o211ai_2
X_10245_ net794 net38 VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__and2_1
X_17841_ _08659_ _08700_ VGND VGND VPWR VPWR _08702_ sky130_fd_sc_hd__nand2_1
XFILLER_121_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17772_ _08563_ _08566_ _08564_ VGND VGND VPWR VPWR _08634_ sky130_fd_sc_hd__o21ai_1
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14984_ _05781_ _05879_ _05880_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__nand3b_1
X_16723_ net620 net1090 net484 net480 VGND VGND VPWR VPWR _07594_ sky130_fd_sc_hd__and4_1
XFILLER_93_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19511_ _00578_ _00699_ _00700_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__nand3_4
X_13935_ net735 net699 VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__nand2_1
X_16654_ net558 net533 net529 net566 VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__a22oi_1
XFILLER_90_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13866_ _04723_ _04726_ _04769_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19442_ _00621_ _00608_ _00607_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__nand3_1
X_15605_ _09199_ _09581_ net1070 _06480_ _06479_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__o221ai_4
XFILLER_90_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12817_ net645 b_h\[9\] VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__nand2_1
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16585_ a_l\[6\] net496 VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__nand2_1
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19373_ _00546_ net230 net621 net717 VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__nand4_2
X_13797_ _02082_ net805 _04607_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15536_ _06414_ _06416_ _06412_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__a21o_1
X_18324_ _09126_ _09127_ _09172_ VGND VGND VPWR VPWR _09173_ sky130_fd_sc_hd__o21ai_2
X_12748_ _03671_ _03674_ _03675_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__nand3_1
X_12679_ net793 _03608_ _03609_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__and3_1
X_18255_ _09101_ _09100_ VGND VGND VPWR VPWR _09102_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_41_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15467_ net223 _06357_ _06324_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__o21a_1
XFILLER_129_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _08063_ _08066_ _08070_ VGND VGND VPWR VPWR _08074_ sky130_fd_sc_hd__a21oi_2
X_18186_ _09025_ _09031_ _09032_ VGND VGND VPWR VPWR _09033_ sky130_fd_sc_hd__nand3_2
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14418_ _05297_ _05298_ _05318_ _05320_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__o2bb2ai_2
X_17137_ _07850_ _07860_ _07851_ VGND VGND VPWR VPWR _08006_ sky130_fd_sc_hd__a21o_1
X_15398_ _06247_ _06248_ _06240_ _06289_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__a31oi_1
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap324 _02876_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_1
Xmax_cap335 _09612_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_4
Xmax_cap313 _05434_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_2
X_14349_ _05249_ _05252_ _05088_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__nand3_1
XFILLER_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap346 _06545_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_1
X_17068_ _07783_ _07792_ _07934_ net343 VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__a22o_1
Xmax_cap357 _03003_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_6
XFILLER_143_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16019_ _06771_ _06775_ _06773_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__a21oi_2
Xmax_cap379 _07530_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_2
XFILLER_66_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19709_ b_l\[9\] net567 VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__nand2_2
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_140_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20415_ clknet_leaf_31_clk _00055_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20346_ net794 net42 VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__and2_2
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20277_ _01519_ _01520_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_147_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11981_ _02882_ _02913_ _02914_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__nand3_4
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10932_ _01878_ _01875_ _01877_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__a21oi_1
XFILLER_44_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13720_ _01888_ _04260_ _04492_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_67_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10863_ net793 net1291 VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__and2_1
X_13651_ _04559_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__inv_2
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10794_ p_hl\[25\] p_lh\[25\] VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__and2_1
X_16370_ net1004 net1023 VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__nand2_1
X_12602_ _03451_ _03528_ _03530_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__nand3_1
X_13582_ _04489_ _04490_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__nand2_1
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12533_ _09417_ _09679_ VGND VGND VPWR VPWR _03465_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15321_ _06214_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__nand2_1
X_18040_ _08888_ _08889_ VGND VGND VPWR VPWR _08890_ sky130_fd_sc_hd__nand2_1
X_15252_ _06072_ _06078_ _06146_ net65 VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__a31o_1
X_12464_ _03394_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__nand2_1
X_14203_ _05084_ _05090_ _05085_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__a21oi_2
X_11415_ _01857_ _02278_ _02274_ _02276_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__o22ai_4
X_12395_ _03324_ _03306_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__nand2_1
X_15183_ _06063_ _06058_ _06056_ _06059_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ _02169_ _02285_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__nand2_1
X_19991_ net735 net551 VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__nand2_4
X_14134_ _04969_ _05035_ _05038_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__nand3_2
XFILLER_140_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18942_ _09796_ _09830_ VGND VGND VPWR VPWR _09834_ sky130_fd_sc_hd__nand2_1
X_14065_ _04884_ _04885_ _04904_ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11277_ _02151_ _02217_ _02218_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__nand3_2
X_13016_ _03942_ VGND VGND VPWR VPWR _03943_ sky130_fd_sc_hd__inv_2
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10228_ net478 VGND VGND VPWR VPWR _09668_ sky130_fd_sc_hd__inv_8
X_18873_ _09745_ _09746_ _09760_ _09761_ VGND VGND VPWR VPWR _09765_ sky130_fd_sc_hd__a22o_1
XFILLER_121_583 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17824_ _08683_ _08674_ _08682_ VGND VGND VPWR VPWR _08685_ sky130_fd_sc_hd__nand3b_2
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17755_ _08617_ VGND VGND VPWR VPWR _08618_ sky130_fd_sc_hd__inv_2
X_14967_ _05793_ _05861_ _05862_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__and3_1
X_16706_ _07433_ _07575_ _07576_ VGND VGND VPWR VPWR _07578_ sky130_fd_sc_hd__nand3_1
XFILLER_63_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17686_ _08526_ _08547_ VGND VGND VPWR VPWR _08549_ sky130_fd_sc_hd__nand2_1
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13918_ _04688_ _04689_ _04690_ _04821_ _04823_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__a32oi_2
X_14898_ net750 net640 VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__nand2_2
X_16637_ _07507_ _07508_ VGND VGND VPWR VPWR _07509_ sky130_fd_sc_hd__nand2_2
X_19425_ _00605_ _00593_ _00604_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__nand3_2
X_13849_ _04750_ _04751_ _04742_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__nand3_4
X_16568_ _07434_ _07435_ _07439_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__nand3_1
X_19356_ _00491_ _00532_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__nand2_1
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15519_ _09581_ _09592_ _06402_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__or3_4
X_18307_ net779 net593 VGND VGND VPWR VPWR _09154_ sky130_fd_sc_hd__nand2_1
X_16499_ net559 net541 VGND VGND VPWR VPWR _07372_ sky130_fd_sc_hd__nand2_1
X_19287_ net760 net755 net575 net567 VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__nand4_4
X_18238_ _09045_ _09082_ _09083_ VGND VGND VPWR VPWR _09085_ sky130_fd_sc_hd__nand3_2
XFILLER_128_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold402 term_low\[4\] VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
X_18169_ _09013_ net305 VGND VGND VPWR VPWR _09017_ sky130_fd_sc_hd__nand2_1
Xhold413 p_hh\[11\] VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 p_hh_pipe\[26\] VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold435 p_ll\[10\] VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
X_20200_ _01440_ net214 VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__nand2_1
XFILLER_145_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap154 _07049_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
Xhold468 p_hh_pipe\[19\] VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap165 _04318_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
Xhold457 p_ll_pipe\[17\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 p_ll_pipe\[26\] VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
X_20131_ net568 net721 VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__and2_1
Xmax_cap198 _04120_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xhold479 p_ll_pipe\[29\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20062_ net735 net549 VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_142_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11200_ _02055_ _02056_ _01991_ _02137_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__o211a_1
X_12180_ _03112_ _03113_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__nand2_1
X_11131_ _02065_ _02070_ _02069_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__o21ai_1
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20329_ net793 net12 VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__and2_1
XFILLER_0_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11062_ net1061 net538 VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__nand2_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15870_ _06745_ _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__nor2_2
XFILLER_95_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14821_ _09308_ _09460_ _05718_ _05719_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__o211ai_2
XFILLER_63_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11964_ net1036 net633 net546 net537 VGND VGND VPWR VPWR _02900_ sky130_fd_sc_hd__nand4_4
X_17540_ _08400_ _08396_ net415 _08401_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__o211ai_4
X_14752_ net163 _05652_ _05538_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__a21bo_1
X_10915_ net713 net707 net441 net364 VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__a31oi_1
X_11895_ _02827_ _02829_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__a21oi_1
X_17471_ _08333_ _08300_ _08332_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__nand3_1
X_13703_ net456 _04609_ net762 net683 VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__o211a_1
X_14683_ net425 _05577_ net426 _05566_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__a31oi_4
X_16422_ _07081_ _07085_ _07289_ _07292_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__nand4_1
X_10846_ net795 net1296 VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__and2_1
XFILLER_71_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13634_ _04538_ _04537_ _04505_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__nand3_4
X_19210_ _10076_ _10102_ _10103_ _10073_ VGND VGND VPWR VPWR _10107_ sky130_fd_sc_hd__a31oi_2
X_16353_ _07095_ _07102_ _07098_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__a21o_1
XFILLER_9_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19141_ _09947_ _09948_ _09937_ VGND VGND VPWR VPWR _10033_ sky130_fd_sc_hd__o21ai_1
X_10777_ p_hl\[23\] p_lh\[23\] VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__and2_1
X_13565_ _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__inv_2
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15304_ _06188_ _06190_ _06196_ _06197_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__o211ai_2
X_16284_ _07157_ _07088_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__nand2_2
X_12516_ net322 _03447_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__nand2_1
X_13496_ _04337_ _04403_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__nand2_1
X_19072_ _09837_ _09793_ VGND VGND VPWR VPWR _09963_ sky130_fd_sc_hd__nand2_1
XFILLER_12_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12447_ _03295_ _03337_ _03339_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__nand3_1
X_18023_ _08870_ _08871_ VGND VGND VPWR VPWR _08873_ sky130_fd_sc_hd__nand2_2
X_15235_ _06047_ _06128_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15166_ _05897_ _06062_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__nor2_1
XFILLER_126_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12378_ net665 net995 VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_93_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14117_ _05019_ _05007_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__nand2_1
X_11329_ _02268_ _02269_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__nand2_1
XFILLER_113_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19974_ _01195_ net589 _01193_ net717 VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__nand4_1
X_15097_ _05992_ _05993_ _09384_ _09449_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_140_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14048_ _04952_ _04953_ _04833_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__a21oi_1
X_18925_ net921 net786 net557 net553 VGND VGND VPWR VPWR _09817_ sky130_fd_sc_hd__nand4_4
X_18856_ _09603_ _09604_ _09609_ VGND VGND VPWR VPWR _09748_ sky130_fd_sc_hd__a21oi_1
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17807_ _08667_ _08668_ VGND VGND VPWR VPWR _08669_ sky130_fd_sc_hd__and2b_1
X_15999_ net607 net515 VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__and2_4
XTAP_TAPCELL_ROW_124_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18787_ _09498_ _09500_ _09502_ VGND VGND VPWR VPWR _09678_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17738_ _09275_ _09679_ _08596_ _08597_ VGND VGND VPWR VPWR _08601_ sky130_fd_sc_hd__o211ai_1
XFILLER_82_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17669_ _08527_ _08528_ _08532_ VGND VGND VPWR VPWR _08533_ sky130_fd_sc_hd__nand3_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19408_ _00470_ _00467_ _00463_ _00468_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_62_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20680_ clknet_leaf_55_clk _00320_ VGND VGND VPWR VPWR p_hl\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19339_ _00512_ _00514_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__nand2_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20114_ _00976_ _00975_ _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__nand3_4
X_20045_ _01179_ _01187_ _01274_ net797 VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__a31o_1
XFILLER_86_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10700_ p_hl\[12\] p_lh\[12\] VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__and2_1
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _02612_ _02614_ _02607_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__a21o_1
X_10631_ p_hl\[1\] p_lh\[1\] p_hl\[0\] net1326 VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__o211ai_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10562_ net794 net1315 VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__and2_1
X_13350_ net714 net751 net1076 net757 VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__a22oi_2
X_12301_ _03220_ _03230_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__nand2_1
X_13281_ net784 net986 VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__nand2_1
X_10493_ _01641_ _01642_ _01650_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__nand3_1
X_12232_ _03164_ _03146_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__nand2_2
X_15020_ _05812_ net310 _05813_ _05673_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__nand4_4
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12163_ _03096_ _03097_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__nor2_1
XFILLER_107_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_75_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _01991_ _01994_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__nor2_1
X_16971_ _07631_ net279 _07778_ _07836_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__o211ai_4
X_12094_ _02991_ _02994_ net293 _03027_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__o211a_1
X_11045_ _01901_ _01938_ _01989_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__nor3_2
X_15922_ _06658_ _06797_ _06791_ _06796_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__o211ai_1
XFILLER_122_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18710_ _09333_ _09465_ _09462_ VGND VGND VPWR VPWR _09594_ sky130_fd_sc_hd__o21a_1
X_19690_ net271 _00893_ _00738_ _00769_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15853_ _06570_ _06644_ VGND VGND VPWR VPWR _06732_ sky130_fd_sc_hd__nand2_1
XFILLER_64_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18641_ _09512_ _09518_ VGND VGND VPWR VPWR _09519_ sky130_fd_sc_hd__nand2_1
XFILLER_18_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15784_ net632 net502 _06659_ _06661_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__a22o_1
X_18572_ _09223_ _09431_ _09429_ _09423_ VGND VGND VPWR VPWR _09443_ sky130_fd_sc_hd__o2bb2ai_1
X_12996_ _03728_ _03919_ _03920_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__nand3b_2
X_14804_ _05702_ _05703_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_24_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11947_ net658 net518 VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__nand2_1
X_17523_ _02589_ _07100_ _08384_ _08386_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__o211a_1
XFILLER_55_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14735_ _05629_ _05632_ _05599_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__a21o_1
XFILLER_17_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11878_ _02435_ _02437_ _02560_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__o21ai_1
X_17454_ _02589_ _06985_ net596 net476 _08318_ VGND VGND VPWR VPWR _08320_ sky130_fd_sc_hd__o2111a_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14666_ _05271_ _05446_ _05441_ _05444_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__o22ai_2
X_16405_ _07274_ _07276_ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__nand2_1
X_17385_ net606 net472 VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__nand2_1
X_10829_ _01842_ _01846_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__nor2_1
XFILLER_60_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13617_ _04417_ _04420_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__nand2_1
X_14597_ _05494_ _05495_ _05496_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_15_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16336_ _07142_ _07138_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__nor2_1
X_13548_ _04434_ _04436_ _04454_ _04455_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_9_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19124_ net760 net575 VGND VGND VPWR VPWR _10014_ sky130_fd_sc_hd__nand2_1
X_16267_ _06957_ _06962_ _06959_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__a21oi_1
X_19055_ _09939_ _09943_ VGND VGND VPWR VPWR _09946_ sky130_fd_sc_hd__nand2_1
X_18006_ _09690_ _08855_ _08856_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__and3_1
X_13479_ _04381_ _04312_ _04252_ _04251_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__and4_4
XPHY_EDGE_ROW_33_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15218_ _06101_ _06105_ _06113_ _06104_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__o211ai_2
X_16198_ _02338_ _06480_ _07066_ _07068_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__o211ai_1
XFILLER_126_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15149_ _06002_ net946 _06042_ _06043_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__o211ai_2
X_19957_ _01176_ _01180_ _01179_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__o21a_1
XFILLER_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18908_ net775 net770 net576 net568 VGND VGND VPWR VPWR _09800_ sky130_fd_sc_hd__and4_1
XFILLER_95_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19888_ _01101_ _01102_ _01098_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__o21ai_1
XFILLER_95_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18839_ _09588_ _09591_ _09580_ _09586_ VGND VGND VPWR VPWR _09732_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_42_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20801_ clknet_leaf_3_clk _00441_ VGND VGND VPWR VPWR b_h\[7\] sky130_fd_sc_hd__dfxtp_4
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20732_ clknet_leaf_35_clk _00372_ VGND VGND VPWR VPWR p_ll\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20663_ clknet_leaf_1_clk _00303_ VGND VGND VPWR VPWR p_hh\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20594_ clknet_leaf_14_clk _00234_ VGND VGND VPWR VPWR p_hh_pipe\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_136_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20028_ _01256_ _01200_ _01254_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__nand3_2
XFILLER_19_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12850_ _03725_ _03774_ _03776_ VGND VGND VPWR VPWR _03779_ sky130_fd_sc_hd__nand3b_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11801_ net637 net537 VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__nand2_2
XFILLER_74_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer91 a_l\[1\] VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd1_1
X_12781_ _03612_ _03697_ _03696_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a21boi_1
Xrebuffer80 b_l\[6\] VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd1_1
X_14520_ net756 net750 net662 net655 VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__nand4_4
XFILLER_27_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11732_ _02665_ _02667_ net227 VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__a21o_1
X_11663_ _02600_ net326 VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__nand2_1
X_14451_ _05351_ _05352_ _05341_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_12_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17170_ _07982_ _08034_ _08033_ net612 net472 VGND VGND VPWR VPWR _08038_ sky130_fd_sc_hd__a32o_1
X_13402_ _04310_ _04311_ _04254_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a21o_1
X_10614_ net794 net1246 VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__and2_1
XFILLER_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14382_ net778 net636 VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__nand2_1
X_16121_ net570 net543 VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__nand2_1
X_11594_ _02528_ _02529_ _02530_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nand3_2
X_13333_ _04217_ _04244_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__nand2_1
X_10545_ net793 net1273 VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_77_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap709 net1076 VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__buf_6
XFILLER_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10476_ _01624_ _01628_ _01631_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__and3_1
X_16052_ _06926_ _06927_ _06853_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__a21boi_1
Xrebuffer181 net977 VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlymetal6s2s_1
X_13264_ _09690_ _04177_ _04178_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__and3_1
Xrebuffer192 _04626_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__buf_2
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12215_ net638 net526 VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__nand2_1
X_13195_ _04113_ _04114_ _04116_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__a21oi_1
X_15003_ _05896_ _05899_ net715 a_h\[6\] VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nand4_1
X_12146_ _03076_ _03074_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__nand2_4
XFILLER_97_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19811_ _09286_ _09308_ _01023_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__o21ai_1
X_16954_ _07113_ _07821_ _07820_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__o21ai_2
X_12077_ net906 net518 _03009_ _03011_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__a22oi_1
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19742_ _00896_ _00947_ _00948_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__nand3_2
X_15905_ _06769_ _06770_ _06778_ _06780_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__o2bb2ai_1
X_11028_ _01964_ _01969_ _01972_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__o21ai_1
X_16885_ net594 net586 net498 net493 VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__nand4_4
XFILLER_77_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19673_ net822 net556 net552 net880 VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__a22oi_1
X_15836_ _06668_ _06669_ _06711_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__o21ai_2
X_18624_ net1131 net589 net581 net775 VGND VGND VPWR VPWR _09500_ sky130_fd_sc_hd__a22oi_1
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15767_ _06645_ _06646_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__nand2_1
XFILLER_64_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18555_ _09419_ _09420_ _09402_ _09403_ VGND VGND VPWR VPWR _09425_ sky130_fd_sc_hd__o211ai_1
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12979_ net1049 net634 net857 net824 VGND VGND VPWR VPWR _03906_ sky130_fd_sc_hd__nand4_4
X_15698_ net628 net632 net512 net505 VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__and4_2
X_17506_ _08360_ _08361_ VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__nand2_1
X_18486_ _09337_ _09342_ _09344_ _09345_ VGND VGND VPWR VPWR _09349_ sky130_fd_sc_hd__o211ai_1
X_14718_ _09308_ _09449_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__o21ai_1
X_17437_ _08171_ _08168_ _08169_ VGND VGND VPWR VPWR _08303_ sky130_fd_sc_hd__a21oi_2
X_14649_ _05464_ _05497_ _05498_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_31_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_27 _09657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_16 _00435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17368_ _08201_ _08202_ _08232_ VGND VGND VPWR VPWR _08235_ sky130_fd_sc_hd__nand3_2
X_19107_ _09996_ _09997_ _09857_ VGND VGND VPWR VPWR _09998_ sky130_fd_sc_hd__a21oi_1
X_16319_ net816 net496 net491 net620 VGND VGND VPWR VPWR _07193_ sky130_fd_sc_hd__a22oi_4
X_17299_ _08104_ _08107_ _08109_ VGND VGND VPWR VPWR _08166_ sky130_fd_sc_hd__o21ai_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput101 net101 VGND VGND VPWR VPWR p[41] sky130_fd_sc_hd__buf_2
XFILLER_134_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19038_ b_l\[2\] net557 VGND VGND VPWR VPWR _09929_ sky130_fd_sc_hd__nand2_1
Xoutput112 net112 VGND VGND VPWR VPWR p[51] sky130_fd_sc_hd__buf_2
Xoutput123 net123 VGND VGND VPWR VPWR p[61] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_132_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_39_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_83_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20715_ clknet_leaf_20_clk _00355_ VGND VGND VPWR VPWR p_lh\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20646_ clknet_leaf_16_clk _00286_ VGND VGND VPWR VPWR p_hh\[12\] sky130_fd_sc_hd__dfxtp_1
Xwire228 _02127_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_2
Xwire239 _06576_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__buf_2
Xwire217 _09706_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__buf_1
Xwire206 _10113_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_4
X_20577_ clknet_leaf_18_clk _00217_ VGND VGND VPWR VPWR p_hh_pipe\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10330_ _00956_ _00967_ _00999_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__o21ai_1
XFILLER_118_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10261_ net794 net1295 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__and2_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12000_ _02934_ _02823_ _02932_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__nand3_2
XFILLER_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ net580 VGND VGND VPWR VPWR _09275_ sky130_fd_sc_hd__inv_8
XFILLER_120_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13951_ _04850_ _04853_ _04838_ _04849_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__o211ai_1
XFILLER_143_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ _09635_ _03826_ _03829_ VGND VGND VPWR VPWR _03830_ sky130_fd_sc_hd__o21ai_1
XFILLER_46_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16670_ net379 _07536_ _07538_ _07520_ VGND VGND VPWR VPWR _07542_ sky130_fd_sc_hd__o211ai_4
XFILLER_62_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13882_ _04779_ _04783_ _04784_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__nand3_1
X_15621_ _06426_ _06456_ _06500_ _06501_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__a2bb2o_1
X_12833_ _03761_ _03677_ _03760_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__nand3_2
XFILLER_27_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15552_ _06433_ _06434_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__or2_1
X_12764_ _03621_ _03623_ _03690_ _03691_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__nand4_2
X_18340_ _09038_ _09042_ _09187_ VGND VGND VPWR VPWR _09191_ sky130_fd_sc_hd__a21o_1
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11715_ _02650_ net507 net682 VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__nand3_1
X_18271_ net804 net759 VGND VGND VPWR VPWR _09117_ sky130_fd_sc_hd__nand2_1
XFILLER_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14503_ _05401_ _05403_ _05264_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__o21ba_1
X_15483_ net716 net640 net635 net719 VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__a22o_1
XFILLER_147_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17222_ _07963_ _07975_ _07965_ VGND VGND VPWR VPWR _08090_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ net674 net481 VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__nand2_1
XFILLER_128_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11646_ _02579_ _02580_ _02578_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__o21ai_1
X_14434_ _01888_ net455 b_l\[14\] net703 _05332_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__o2111ai_4
XFILLER_11_860 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17153_ _08017_ _08019_ _08021_ VGND VGND VPWR VPWR _08022_ sky130_fd_sc_hd__o21a_1
X_11577_ _02487_ _02488_ net359 _02512_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__nand4_1
XFILLER_7_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput25 a[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 b[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 a[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xwire740 net742 VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__buf_12
X_14365_ _05183_ _05185_ _05190_ _05237_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__a22oi_4
X_10528_ net1311 _01673_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__nor2_1
XFILLER_128_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16104_ net572 net541 VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__nand2_1
X_17084_ net582 net498 VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__nand2_1
Xmax_cap506 net509 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__buf_6
X_13316_ _04223_ _04225_ _04220_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a21o_1
X_14296_ _05053_ _05054_ _05052_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__a21oi_1
Xinput47 b[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 b[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
X_16035_ _06907_ _06796_ _06908_ _06910_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__nand4_4
Xmax_cap528 net529 VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_12
Xmax_cap539 b_h\[1\] VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__buf_8
X_13247_ net787 net693 VGND VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand2_1
X_10459_ _01620_ _01621_ _01622_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_114_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13178_ _04099_ _09668_ net634 VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__or3b_1
X_12129_ _03045_ _03046_ _03063_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__o21ai_2
X_17986_ net623 net779 VGND VGND VPWR VPWR _08837_ sky130_fd_sc_hd__nand2_2
XFILLER_111_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16937_ net344 _07636_ _07655_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__a21boi_1
X_19725_ _00927_ _00931_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__nand2_1
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16868_ net612 net479 VGND VGND VPWR VPWR _07738_ sky130_fd_sc_hd__nand2_1
XFILLER_92_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19656_ _00853_ _00854_ _00856_ _00857_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__a31oi_1
XFILLER_38_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15819_ _06696_ _06697_ _09188_ _09602_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__o2bb2a_1
X_16799_ _07498_ _07668_ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__nand2_2
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18607_ net782 net564 VGND VGND VPWR VPWR _09481_ sky130_fd_sc_hd__nand2_2
X_19587_ _00661_ net408 _00662_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__a21boi_2
X_18538_ net621 net743 net737 net626 VGND VGND VPWR VPWR _09407_ sky130_fd_sc_hd__a22oi_1
XFILLER_80_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20500_ clknet_leaf_16_clk _00140_ VGND VGND VPWR VPWR term_mid\[44\] sky130_fd_sc_hd__dfxtp_1
X_18469_ net610 net754 VGND VGND VPWR VPWR _09331_ sky130_fd_sc_hd__nand2_1
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20431_ clknet_leaf_16_clk _00071_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfxtp_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20362_ clknet_leaf_50_clk _00002_ VGND VGND VPWR VPWR b_l\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_146_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20293_ _01512_ _01518_ _01537_ _01538_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__a211oi_1
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_145_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11500_ _02436_ _02434_ _02433_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__nand3_1
XFILLER_51_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12480_ _03406_ _03408_ _03270_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_22_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _02366_ _02355_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__nand2_2
X_20629_ clknet_leaf_49_clk _00269_ VGND VGND VPWR VPWR p_ll_pipe\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ _02290_ net360 VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__nand2_1
X_14150_ _05053_ _05054_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__nand2_2
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13101_ _03981_ _03985_ _04024_ _04025_ VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__a22o_1
X_10313_ term_low\[24\] term_mid\[24\] VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__xor2_1
X_11293_ _02149_ _02228_ _02229_ _02141_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__a31oi_4
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081_ _04983_ _04984_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__nand2_2
XFILLER_133_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13032_ _03901_ _03913_ _03916_ VGND VGND VPWR VPWR _03958_ sky130_fd_sc_hd__o21ai_4
X_10244_ net794 net37 VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__and2_1
X_17840_ _08658_ _08697_ _08699_ _08655_ VGND VGND VPWR VPWR _08701_ sky130_fd_sc_hd__nand4_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17771_ _08631_ net477 net899 _08630_ VGND VGND VPWR VPWR _08633_ sky130_fd_sc_hd__nand4_4
XFILLER_75_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19510_ _00697_ _00695_ _00696_ _00577_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__o211ai_4
X_14983_ _05877_ _05878_ _05781_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__a21oi_4
X_16722_ net1090 net484 net480 net620 VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__a22o_1
X_13934_ _04779_ _04782_ _04784_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__o21ai_1
X_16653_ net559 net533 VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13865_ _04725_ _04718_ _04724_ _04766_ _04767_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__o2111ai_1
X_19441_ _00607_ _00608_ _00617_ _00618_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15604_ _06475_ _06481_ VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__nand2_1
X_12816_ net648 b_h\[10\] VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__nand2_1
XFILLER_62_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19372_ _00546_ net230 _00545_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__and3_1
X_16584_ net928 net491 VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__nand2_1
X_18323_ _09170_ _09171_ VGND VGND VPWR VPWR _09172_ sky130_fd_sc_hd__nand2_1
X_13796_ _09220_ _09439_ _02082_ net922 VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__o22a_1
XFILLER_97_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15535_ _06414_ _06416_ _06412_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__a21oi_1
X_12747_ _03671_ _03674_ _03675_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__and3_1
XFILLER_147_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12678_ _03605_ net136 _03602_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__a21o_1
X_18254_ _09021_ _08951_ _09020_ VGND VGND VPWR VPWR _09101_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_41_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15466_ _06356_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__inv_2
X_11629_ _02441_ _02567_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_116_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _08047_ _08050_ _08071_ _08072_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__o211ai_2
X_18185_ _09026_ net759 net623 VGND VGND VPWR VPWR _09032_ sky130_fd_sc_hd__nand3_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14417_ _05300_ _05307_ _05309_ _05314_ _05312_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__o311a_1
XFILLER_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_129_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17136_ _07998_ _08000_ _07895_ VGND VGND VPWR VPWR _08005_ sky130_fd_sc_hd__o21ai_1
X_15397_ _06283_ _06287_ _06286_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap314 _05174_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__buf_6
X_14348_ _05251_ _05106_ _05250_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__nand3_4
XFILLER_143_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap358 _02872_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_4
X_17067_ _07782_ _07791_ _07934_ net343 VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__a2bb2oi_2
Xmax_cap369 _09879_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_2
X_14279_ net315 _05141_ _05182_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__o21ai_2
Xmax_cap347 _06103_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_2
X_16018_ _06771_ _06775_ _06773_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__a21o_1
XFILLER_97_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17969_ net623 net790 net781 net615 VGND VGND VPWR VPWR _08821_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_127_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19708_ net574 b_l\[10\] VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__nand2_1
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19639_ _00726_ _00728_ _00835_ _00836_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__a22o_1
XFILLER_92_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20414_ clknet_leaf_30_clk _00054_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20345_ net794 net41 VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_8_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20276_ _01519_ _01520_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__nand2_1
XFILLER_103_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11980_ _02744_ _02881_ _02911_ _02912_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__o211ai_4
XFILLER_91_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10931_ _01876_ _01866_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__nand2_1
XFILLER_84_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10862_ net793 net1249 VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__and2_1
X_13650_ _04438_ net352 _04451_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__a21bo_1
X_10793_ p_hl\[25\] p_lh\[25\] VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nor2_1
X_12601_ _03528_ _03530_ _03425_ _03448_ VGND VGND VPWR VPWR _03532_ sky130_fd_sc_hd__o2bb2ai_2
X_13581_ net757 net694 VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__nand2_2
XFILLER_24_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12532_ _03380_ _03458_ _03459_ VGND VGND VPWR VPWR _03464_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_80_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15320_ _06075_ _06212_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__nand2_2
X_12463_ net437 _03391_ _03393_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__nand3_4
X_15251_ _06072_ _06078_ _06146_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__a21oi_1
X_11414_ _02351_ _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__nor2_1
XFILLER_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14202_ _05086_ _05092_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__nand2_1
XFILLER_138_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12394_ _03304_ _03305_ _03321_ _03323_ VGND VGND VPWR VPWR _03327_ sky130_fd_sc_hd__o211ai_2
X_15182_ net65 _06077_ _06078_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__nor3b_1
X_11345_ _02165_ _02168_ _02171_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__o21ai_1
XFILLER_4_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19990_ net731 net563 VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__nand2_1
X_14133_ _05004_ _05006_ _05025_ _05029_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__o2bb2ai_1
X_11276_ _02185_ _02186_ _02203_ _02206_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_111_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18941_ _09824_ _09826_ _09807_ VGND VGND VPWR VPWR _09833_ sky130_fd_sc_hd__a21o_1
XFILLER_4_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14064_ _04914_ _04908_ _04913_ _04939_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__a22oi_2
X_10227_ net486 VGND VGND VPWR VPWR _09657_ sky130_fd_sc_hd__inv_6
X_13015_ _03799_ _03941_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__nand2_1
XFILLER_4_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18872_ net411 _09746_ _09760_ _09761_ VGND VGND VPWR VPWR _09764_ sky130_fd_sc_hd__nand4_2
XFILLER_121_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17823_ _09646_ _08673_ _08681_ _08683_ VGND VGND VPWR VPWR _08684_ sky130_fd_sc_hd__o22ai_2
X_17754_ _08457_ _08542_ _08541_ VGND VGND VPWR VPWR _08617_ sky130_fd_sc_hd__a21boi_2
X_14966_ _05861_ _05862_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nand2_1
X_16705_ _07575_ _07576_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__nand2_1
X_13917_ _04821_ _04823_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__nand2_1
XFILLER_48_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17685_ _08478_ _08525_ _08524_ VGND VGND VPWR VPWR _08548_ sky130_fd_sc_hd__o21ai_1
X_19424_ _00602_ _00598_ _00594_ _00603_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__o211ai_4
X_14897_ _05794_ _05795_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__nand2_2
X_16636_ net453 _07502_ _07506_ _07492_ VGND VGND VPWR VPWR _07508_ sky130_fd_sc_hd__o211ai_4
X_13848_ _04750_ _04751_ _04742_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__a21oi_1
X_16567_ _07434_ _07435_ _07184_ _07307_ net145 VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__a221o_1
XFILLER_95_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13779_ _04585_ _04683_ _04685_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__nand3_2
XFILLER_16_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19355_ _00528_ _00529_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__nand2_1
X_15518_ net1105 net540 net848 _06403_ net797 VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__a311oi_1
X_18306_ _09155_ _09242_ VGND VGND VPWR VPWR _09153_ sky130_fd_sc_hd__nor2_1
X_19286_ net575 net567 net458 VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__and3_1
X_16498_ _09340_ _09581_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__nor2_1
X_18237_ _09082_ _09083_ VGND VGND VPWR VPWR _09084_ sky130_fd_sc_hd__nand2_1
X_15449_ _06214_ _06215_ _06339_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__a21oi_4
XFILLER_117_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18168_ _08895_ _08896_ _09003_ _09010_ net1118 VGND VGND VPWR VPWR _09016_ sky130_fd_sc_hd__o221ai_4
XFILLER_144_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold425 mid_sum\[26\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 p_hh\[10\] VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 p_hh_pipe\[27\] VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap144 _07719_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
X_17119_ _07986_ _07987_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__nand2_1
Xhold403 p_ll_pipe\[7\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ _08939_ _08945_ _08941_ VGND VGND VPWR VPWR _08948_ sky130_fd_sc_hd__nor3_4
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold458 mid_sum\[22\] VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 p_hh\[17\] VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap177 _03084_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_2
XFILLER_89_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20130_ _01297_ _01293_ _01295_ _01365_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__o211ai_4
Xhold447 p_ll_pipe\[21\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap199 _03098_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
XFILLER_98_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap188 net189 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20061_ net731 net557 VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__nand2_1
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11130_ _02071_ _02072_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__nand2_1
X_20328_ net793 net1 VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__and2_1
XFILLER_134_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_79_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11061_ net678 net965 net538 net681 VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20259_ _01462_ _01463_ _01466_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__a21o_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14820_ _05718_ _05719_ _05715_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__a21o_1
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11963_ net633 net537 VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__nand2_4
X_14751_ _05650_ _05642_ _05540_ _05651_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__o211ai_4
X_11894_ net708 net475 _02827_ _02828_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__a22oi_1
X_10914_ _01859_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__xnor2_1
X_17470_ _08333_ _08300_ _08332_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__and3_1
XFILLER_60_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13702_ net924 net768 net676 net673 VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__nand4_1
X_14682_ _05576_ _05577_ net426 VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__nand3_4
XFILLER_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16421_ _07293_ _07294_ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__nand2_1
X_10845_ net795 net1164 VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_88_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13633_ _04505_ _04538_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__nand2_4
X_16352_ _07108_ _07119_ _07109_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__a21boi_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19140_ _10030_ _10031_ VGND VGND VPWR VPWR _10032_ sky130_fd_sc_hd__nand2_2
X_10776_ p_hl\[23\] p_lh\[23\] VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__nor2_1
X_13564_ _04465_ _04467_ _04471_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__nand3_4
X_15303_ _06196_ _06197_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__nand2_1
X_16283_ _07156_ _07087_ _07155_ _07086_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__nand4_4
X_12515_ _03262_ _03441_ _03440_ net354 VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__o211ai_4
X_13495_ net768 net689 net683 net924 VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__a22oi_2
X_19071_ _09958_ _09959_ _09924_ VGND VGND VPWR VPWR _09962_ sky130_fd_sc_hd__a21o_1
X_12446_ _03298_ _03334_ _03335_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__nand3_1
X_18022_ net781 net886 net605 net790 VGND VGND VPWR VPWR _08872_ sky130_fd_sc_hd__a22oi_2
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15234_ _06047_ _06126_ _06127_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__nand3b_4
X_12377_ net1048 net495 VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15165_ _09384_ _09439_ _05899_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__o21a_1
XFILLER_125_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11328_ _02192_ _02197_ _02263_ _02264_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__nand4_2
XPHY_EDGE_ROW_97_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14116_ _05017_ _05018_ _05009_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__nand3_2
X_19973_ _01193_ net717 net589 VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__nand3_2
X_15096_ _05940_ _05941_ _05948_ _05955_ _05959_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__o2111ai_4
XFILLER_140_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11259_ _09177_ _09613_ _02108_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__o21a_1
XFILLER_113_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14047_ _04950_ _04951_ _04834_ VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__nand3_4
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18924_ net817 net553 VGND VGND VPWR VPWR _09816_ sky130_fd_sc_hd__nand2_2
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18855_ _09745_ _09746_ VGND VGND VPWR VPWR _09747_ sky130_fd_sc_hd__nand2_1
Xsplit153 a_l\[7\] VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__clkbuf_4
X_17806_ _08666_ _08665_ _08664_ VGND VGND VPWR VPWR _08668_ sky130_fd_sc_hd__nand3_1
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15998_ _06860_ _06870_ _06871_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__nand3_4
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18786_ _09638_ _09671_ _09672_ VGND VGND VPWR VPWR _09677_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_124_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17737_ _08596_ _08597_ _08594_ VGND VGND VPWR VPWR _08600_ sky130_fd_sc_hd__a21o_1
XFILLER_48_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14949_ _05692_ _05696_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__nand2_1
X_17668_ _08442_ _08431_ _08429_ VGND VGND VPWR VPWR _08532_ sky130_fd_sc_hd__a21boi_1
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16619_ _07367_ _07408_ net255 VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__a21oi_4
X_19407_ _00505_ _00518_ _00507_ _00516_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__a2bb2o_2
X_17599_ _08458_ _08462_ net795 VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_18_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19338_ _00511_ _00513_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_139_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19269_ net776 net808 net556 net552 VGND VGND VPWR VPWR _10171_ sky130_fd_sc_hd__nand4_2
XFILLER_117_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20113_ _01272_ _01179_ _01269_ _01347_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__o211a_1
X_20044_ _01179_ _01187_ _01274_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__a21oi_1
XFILLER_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10630_ p_hl\[1\] p_lh\[1\] VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__nor2_1
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10561_ net794 net1308 VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__and2_1
X_10492_ term_mid\[48\] term_high\[48\] term_high\[49\] term_high\[50\] term_high\[51\]
+ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__o2111a_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12300_ _03218_ _03219_ _03231_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__nand3_1
XFILLER_108_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13280_ net784 net693 net986 net787 VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__a22o_1
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12231_ _03144_ _03145_ _03162_ _03163_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__nand4_4
Xrebuffer352 b_h\[12\] VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12162_ _03094_ _03095_ net983 net474 VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__and4_1
XFILLER_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11113_ _02055_ _02056_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__nor2_1
XFILLER_123_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16970_ _07835_ _07836_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__nand2_1
X_12093_ _02991_ net294 _03027_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__o21ai_4
XFILLER_77_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _01934_ _01937_ _01987_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__a22oi_2
X_15921_ _06792_ _06798_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__nand2_1
XFILLER_103_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18640_ _09475_ _09513_ _09516_ VGND VGND VPWR VPWR _09518_ sky130_fd_sc_hd__nand3_1
X_15852_ _06643_ _06569_ VGND VGND VPWR VPWR _06731_ sky130_fd_sc_hd__nand2_1
XFILLER_77_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15783_ _06659_ _06661_ net632 net502 VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__nand4_2
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18571_ _09322_ _09440_ _09442_ net794 VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__o211a_1
X_12995_ _03917_ _03918_ _03728_ VGND VGND VPWR VPWR _03922_ sky130_fd_sc_hd__a21oi_1
X_14803_ _05677_ _05699_ _05700_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__nand3b_2
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11946_ _02730_ _02746_ _02744_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__a21oi_2
X_17522_ net1093 net485 _08385_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__a21o_1
X_14734_ _05629_ _05632_ _05599_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__a21oi_1
X_17453_ _02589_ _06985_ _08318_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__o21ai_1
X_11877_ _02812_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nor2_1
X_16404_ _07259_ _07270_ _07272_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__and3_1
XFILLER_72_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _05418_ _05422_ _05421_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__a21boi_2
XFILLER_33_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17384_ _09210_ _09679_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__nor2_1
X_10828_ _01837_ _01843_ _01845_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__a21oi_1
X_13616_ _04521_ _04522_ net777 net673 VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__nand4_1
X_14596_ net349 _05358_ _05494_ _05495_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_15_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16335_ _07199_ _07202_ _07205_ VGND VGND VPWR VPWR _07209_ sky130_fd_sc_hd__nand3_1
X_10759_ _01782_ _01784_ net442 VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__o21a_1
X_13547_ _04434_ _04436_ _04456_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__nand3_2
X_19123_ net589 net749 VGND VGND VPWR VPWR _10013_ sky130_fd_sc_hd__nand2_2
X_16266_ _09188_ _09613_ _06959_ _06961_ _06898_ VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__o32a_1
X_19054_ _09941_ _09943_ net764 net575 VGND VGND VPWR VPWR _09945_ sky130_fd_sc_hd__and4_1
X_18005_ _08851_ _08853_ net338 _08829_ VGND VGND VPWR VPWR _08856_ sky130_fd_sc_hd__nand4b_2
X_13478_ net196 _04381_ _04313_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__nand3_1
X_15217_ _06111_ _06112_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__nor2_2
X_16197_ _07067_ _07069_ net629 net1032 VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__o211ai_1
X_12429_ _03357_ _03360_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__a21o_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15148_ _06037_ _06040_ _06006_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__a21o_1
XFILLER_114_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19956_ _01175_ _01167_ _01085_ _01173_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__o211ai_2
X_15079_ _05971_ _05976_ _05975_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__o21ai_1
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18907_ net770 net576 net568 net775 VGND VGND VPWR VPWR _09799_ sky130_fd_sc_hd__a22oi_1
X_19887_ _00984_ _00987_ _01101_ _01102_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__a211o_1
XFILLER_95_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18838_ _09725_ _09729_ _09728_ VGND VGND VPWR VPWR _09731_ sky130_fd_sc_hd__a21oi_2
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18769_ net1064 net1084 net560 net792 VGND VGND VPWR VPWR _09659_ sky130_fd_sc_hd__a22oi_2
X_20800_ clknet_leaf_3_clk _00440_ VGND VGND VPWR VPWR b_h\[6\] sky130_fd_sc_hd__dfxtp_4
Xclkbuf_leaf_47_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_104_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20731_ clknet_leaf_35_clk _00371_ VGND VGND VPWR VPWR p_ll\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20662_ clknet_leaf_1_clk _00302_ VGND VGND VPWR VPWR p_hh\[28\] sky130_fd_sc_hd__dfxtp_1
X_20593_ clknet_leaf_14_clk _00233_ VGND VGND VPWR VPWR p_hh_pipe\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_137_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_57_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20027_ _01153_ _01253_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__nand2_1
XFILLER_100_384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11800_ _02734_ _02735_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_38_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_8
X_12780_ _03696_ _03708_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__nand2_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer70 a_h\[8\] VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_15_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer81 b_l\[6\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd1_1
X_11731_ _02667_ _02665_ net227 VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__a21oi_4
Xrebuffer92 net888 VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlymetal6s2s_1
X_11662_ _02596_ _02597_ _02575_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__nand3_4
X_14450_ _05349_ _05345_ _05342_ _05350_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_12_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11593_ _02529_ _02528_ _02530_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__a21o_1
X_13401_ _04254_ _04310_ _04311_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__nand3_1
X_10613_ net794 net1201 VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__and2_1
X_14381_ _05162_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__nand2_1
X_10544_ net793 net1258 VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__and2_1
XFILLER_128_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16120_ net595 net521 VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__nand2_1
X_13332_ _04200_ _04216_ _04242_ _04243_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__a22oi_1
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10475_ _01634_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__nor2_1
X_16051_ _06926_ _06927_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__nand2_1
Xrebuffer171 _02804_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__buf_1
Xrebuffer182 _02606_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__buf_2
X_13263_ _04156_ _04176_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__or2_1
Xrebuffer160 net956 VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__buf_6
Xrebuffer193 _02042_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12214_ net647 net518 VGND VGND VPWR VPWR _03148_ sky130_fd_sc_hd__nand2_1
X_13194_ net793 _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__nand2_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15002_ net715 a_h\[6\] _05896_ _05899_ VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__a22o_1
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12145_ _03077_ _03079_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__nand2_1
XFILLER_97_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19810_ _00915_ _01020_ _01015_ _01019_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__o211ai_2
X_16953_ _07819_ _07822_ VGND VGND VPWR VPWR _07823_ sky130_fd_sc_hd__nor2_1
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12076_ _02887_ _03008_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__nand2_2
X_19741_ _00894_ _00895_ _00944_ _00945_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__nand4_2
X_15904_ _06776_ _06777_ _06769_ _06770_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__o211ai_1
X_11027_ _01968_ _01956_ _01967_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__nand3_1
X_16884_ net586 net493 VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__nand2_1
X_19672_ net877 net819 net556 net553 VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__nand4_2
X_15835_ _06709_ _06710_ _06672_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__nand3_1
XFILLER_92_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18623_ net775 net581 VGND VGND VPWR VPWR _09499_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
X_18554_ _09402_ _09403_ _09421_ VGND VGND VPWR VPWR _09424_ sky130_fd_sc_hd__a21o_1
X_15766_ _06567_ _06572_ _06570_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__o21a_1
X_17505_ net796 _08369_ _08370_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__nor3_1
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12978_ net634 net857 VGND VGND VPWR VPWR _03905_ sky130_fd_sc_hd__nand2_1
XFILLER_45_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15697_ net628 net505 VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__nand2_1
X_11929_ net672 net665 net511 net508 VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__nand4_2
XFILLER_72_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18485_ _09343_ _09344_ _09345_ VGND VGND VPWR VPWR _09348_ sky130_fd_sc_hd__a21o_1
X_14717_ _05613_ _05614_ _05616_ _05479_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__o2bb2ai_1
X_17436_ _08168_ _08171_ _08169_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__a21o_1
X_14648_ _05546_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_17 _00436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17367_ _08199_ _08200_ _08232_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__a21boi_1
XANTENNA_28 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16318_ net812 net496 VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19106_ _09625_ _09629_ _09596_ _09991_ _09995_ VGND VGND VPWR VPWR _09997_ sky130_fd_sc_hd__o2111ai_2
X_14579_ net740 net736 net677 net670 VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__nand4_2
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17298_ _07992_ _08134_ _08137_ _08139_ _08040_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__a32o_1
XFILLER_146_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16249_ _07108_ _07109_ _07120_ VGND VGND VPWR VPWR _07124_ sky130_fd_sc_hd__nand3_1
X_19037_ _09811_ _09817_ _09814_ VGND VGND VPWR VPWR _09928_ sky130_fd_sc_hd__a21oi_1
Xoutput102 net102 VGND VGND VPWR VPWR p[42] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR p[52] sky130_fd_sc_hd__buf_2
Xoutput124 net124 VGND VGND VPWR VPWR p[62] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_132_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19939_ _01097_ _01157_ _01158_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__nand3_1
XFILLER_101_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20714_ clknet_leaf_25_clk _00354_ VGND VGND VPWR VPWR p_lh\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20645_ clknet_leaf_16_clk _00285_ VGND VGND VPWR VPWR p_hh\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_23_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire229 _00185_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
X_20576_ clknet_leaf_27_clk _00216_ VGND VGND VPWR VPWR p_hh_pipe\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10260_ net794 net1197 VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__and2_1
XFILLER_127_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ net747 VGND VGND VPWR VPWR _09264_ sky130_fd_sc_hd__inv_16
XFILLER_105_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13950_ _04839_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nand2_1
XFILLER_86_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12901_ _03824_ _03825_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__nand2_2
X_15620_ _06500_ _06501_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__nand2_1
XFILLER_47_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13881_ _04785_ _04786_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_87_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _03739_ _03740_ _03757_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15551_ _09199_ _09526_ _06432_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__o21a_1
X_12763_ _03690_ _03691_ _03624_ VGND VGND VPWR VPWR _03693_ sky130_fd_sc_hd__a21o_1
XFILLER_54_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11714_ _02524_ _02650_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__nand2_1
XFILLER_70_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18270_ net622 net754 VGND VGND VPWR VPWR _09116_ sky130_fd_sc_hd__nand2_1
X_14502_ _05399_ _05400_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__nand2_1
X_15482_ _09362_ _06371_ net635 VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__or3b_1
X_17221_ net451 _07970_ _07973_ _07963_ VGND VGND VPWR VPWR _08089_ sky130_fd_sc_hd__o211a_1
X_12694_ _03621_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__nand2_1
X_14433_ _05332_ _05335_ _05334_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__and3_1
X_11645_ net698 net692 net975 net492 _02578_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__a41o_1
Xinput26 a[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
X_17152_ _07867_ _07885_ _08015_ _08016_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__o211ai_2
X_11576_ _02513_ _02491_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__nand2_2
Xwire730 b_l\[11\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__buf_6
Xinput37 b[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 a[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ _05116_ _05245_ _05239_ _05241_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__o2bb2ai_2
X_10527_ net1371 net1323 net1310 _01669_ net65 VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__a41o_1
X_16103_ _06440_ _06867_ _06861_ _06864_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__o22a_1
Xmax_cap507 net508 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__buf_12
X_17083_ net593 net488 VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__nand2_1
X_13315_ _09155_ _09417_ _04223_ _04225_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__o211ai_1
Xinput48 b[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput59 b[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_14295_ _05195_ _05197_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__nand2_1
X_10458_ _01621_ _01620_ net796 VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__a21oi_1
X_16034_ _06907_ _06908_ _06909_ _06795_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__o2bb2ai_2
Xmax_cap529 net530 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_12
X_13246_ net777 net704 VGND VGND VPWR VPWR _04161_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_114_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10389_ term_mid\[34\] term_high\[34\] _01560_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__a21o_1
XFILLER_124_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13177_ b_h\[15\] _04002_ _04098_ net999 VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__o22a_1
X_12128_ _03061_ _03062_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__nand2_1
XFILLER_111_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17985_ _08819_ net779 net627 _08820_ VGND VGND VPWR VPWR _08836_ sky130_fd_sc_hd__a31o_1
XFILLER_2_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12059_ _02987_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__nor2_1
X_16936_ _07649_ _07650_ _07637_ _07636_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__a31o_1
XFILLER_96_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19724_ _00929_ _00923_ _00928_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__nand3_2
XFILLER_93_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16867_ _07678_ _07683_ _07680_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__a21oi_1
XFILLER_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19655_ _00708_ _00716_ _00855_ net797 VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__a31o_1
X_15818_ net613 net1117 net542 net521 VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__nand4_4
X_16798_ net572 net513 net506 net1069 VGND VGND VPWR VPWR _07669_ sky130_fd_sc_hd__a22oi_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18606_ _09478_ _09479_ VGND VGND VPWR VPWR _09480_ sky130_fd_sc_hd__nand2_2
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19586_ net833 _00781_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__nand2_1
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15749_ _06620_ _06625_ _06624_ _06584_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__o211ai_1
XFILLER_92_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18537_ net621 net626 net743 net737 VGND VGND VPWR VPWR _09405_ sky130_fd_sc_hd__nand4_2
X_18468_ net619 net749 VGND VGND VPWR VPWR _09330_ sky130_fd_sc_hd__nand2_1
XFILLER_33_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17419_ _08230_ _08235_ VGND VGND VPWR VPWR _08285_ sky130_fd_sc_hd__nand2_1
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18399_ _09250_ _09251_ net604 net764 VGND VGND VPWR VPWR _09255_ sky130_fd_sc_hd__and4_1
X_20430_ clknet_leaf_15_clk _00070_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfxtp_1
XFILLER_146_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20361_ clknet_leaf_51_clk _00001_ VGND VGND VPWR VPWR b_l\[1\] sky130_fd_sc_hd__dfxtp_4
X_20292_ _01537_ net168 _01512_ _01518_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__o211a_1
XFILLER_142_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11430_ _02276_ _02283_ net400 _02367_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__o22ai_4
X_20628_ clknet_leaf_47_clk _00268_ VGND VGND VPWR VPWR p_ll_pipe\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20559_ clknet_leaf_18_clk _00199_ VGND VGND VPWR VPWR mid_sum\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11361_ _02298_ _02300_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__nand2_1
XFILLER_4_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13100_ _03976_ _03983_ _03984_ _04023_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__a31o_1
XFILLER_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10312_ _00773_ net1351 _00795_ _00806_ net797 VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__a311oi_1
X_11292_ _02140_ _02131_ _02232_ _02231_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__a22oi_4
XPHY_EDGE_ROW_60_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14080_ net783 net643 net639 net788 VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a22oi_1
XFILLER_79_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13031_ _09471_ _09679_ _03883_ _03881_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__o31a_1
X_10243_ net794 net36 VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__and2_1
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17770_ a_l\[11\] net477 _08630_ _08631_ VGND VGND VPWR VPWR _08632_ sky130_fd_sc_hd__a22o_1
XFILLER_67_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16721_ _07492_ _07506_ net453 _07502_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_59_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14982_ _05770_ _05773_ _05877_ _05878_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__nand4_2
X_13933_ net724 net709 net431 _04836_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__a31o_1
X_16652_ net874 net903 VGND VGND VPWR VPWR _07524_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13864_ _04766_ _04767_ _04727_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__a21o_1
X_19440_ _00617_ _00618_ _00607_ _00608_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__o211ai_2
X_16583_ net812 net1032 VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__nand2_1
X_15603_ _06479_ _06481_ _06475_ VGND VGND VPWR VPWR _06485_ sky130_fd_sc_hd__a21o_1
X_12815_ net654 net490 VGND VGND VPWR VPWR _03744_ sky130_fd_sc_hd__nand2_1
X_19371_ net621 net717 net230 _00546_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__a22o_1
X_15534_ _09144_ _09581_ _06414_ _06416_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__o211ai_1
X_18322_ _09167_ _09132_ _09168_ VGND VGND VPWR VPWR _09171_ sky130_fd_sc_hd__nand3_4
X_13795_ _04655_ _04677_ _04657_ _04659_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__o2bb2ai_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_12746_ _03674_ _03675_ _03671_ VGND VGND VPWR VPWR _03676_ sky130_fd_sc_hd__a21o_1
XFILLER_43_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12677_ _03602_ _03605_ net136 VGND VGND VPWR VPWR _03608_ sky130_fd_sc_hd__nand3_1
X_18253_ _09097_ _09099_ VGND VGND VPWR VPWR _09100_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_41_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15465_ _06347_ _06348_ _06353_ _06354_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__o22ai_1
X_11628_ _02331_ _02438_ _02334_ _02332_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_116_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _08068_ _08070_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__nand2_1
X_18184_ _09027_ net754 net626 VGND VGND VPWR VPWR _09031_ sky130_fd_sc_hd__nand3_1
X_15396_ _06283_ _06287_ _06286_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__o21a_1
X_14416_ _05127_ _05132_ _05313_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17135_ _07896_ _07997_ _08003_ VGND VGND VPWR VPWR _08004_ sky130_fd_sc_hd__o21ai_2
X_14347_ _05246_ _05116_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__nand2_1
XFILLER_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11559_ net652 net537 VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__nand2_1
Xmax_cap315 _05139_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_1
XFILLER_144_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap359 _02510_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_6
X_17066_ _07244_ _07632_ _07931_ _07932_ VGND VGND VPWR VPWR _07935_ sky130_fd_sc_hd__o211ai_2
Xmax_cap337 _08961_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_1
X_14278_ _05177_ _05178_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__nand2_2
Xmax_cap348 _06003_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_6
X_16017_ _06768_ _06856_ _06891_ _06892_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__o211ai_4
XFILLER_124_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13229_ _04138_ net713 net777 _04136_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__a31o_1
XFILLER_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17968_ net623 net790 net781 net615 VGND VGND VPWR VPWR _08820_ sky130_fd_sc_hd__and4_1
XFILLER_69_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_108_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16919_ _07787_ _07788_ VGND VGND VPWR VPWR _07789_ sky130_fd_sc_hd__nand2_1
XFILLER_93_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17899_ net254 _08754_ _08755_ _08756_ VGND VGND VPWR VPWR _08758_ sky130_fd_sc_hd__and4bb_1
XFILLER_84_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19707_ net580 b_l\[11\] VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__nand2_1
XFILLER_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19638_ _00835_ _00836_ _00729_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__a21o_1
XFILLER_38_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19569_ _09264_ _09286_ _00651_ _00653_ _00455_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__o32ai_4
XPHY_EDGE_ROW_117_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20413_ clknet_leaf_30_clk _00053_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfxtp_1
XFILLER_135_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20344_ net794 net40 VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_8_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20275_ _01520_ _01519_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__and2b_1
XFILLER_115_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_126_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10930_ _01876_ net530 net713 VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__and3_1
XFILLER_90_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10861_ net793 net1271 VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__and2_1
X_12600_ _03529_ _03526_ _03527_ _03522_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__a22o_1
XFILLER_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10792_ _01806_ _01807_ _01814_ _01815_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__o31a_1
XFILLER_71_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13580_ net751 net701 VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_135_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12531_ _03381_ _03460_ _03461_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_80_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12462_ _03312_ _03318_ _03390_ _03392_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__o22ai_4
XFILLER_12_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15250_ _06144_ _06145_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__nand2_1
X_11413_ net401 _02347_ _02349_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__a21oi_1
X_14201_ _09690_ _05104_ _05105_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__and3_1
X_12393_ _03306_ _03321_ _03323_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__nand3_1
X_15181_ _06074_ _06076_ _06073_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__o21bai_1
XFILLER_125_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11344_ _02165_ _02171_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__nand2_1
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14132_ _04968_ _05031_ net244 VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__nand3_2
XFILLER_140_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11275_ _02185_ _02186_ _02204_ _02207_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_111_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18940_ _09826_ _09807_ _09824_ VGND VGND VPWR VPWR _09832_ sky130_fd_sc_hd__and3_1
X_14063_ _04913_ _04939_ _04915_ _04909_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__o2bb2ai_2
X_13014_ _03762_ _03768_ _03797_ _03801_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__a31o_1
X_10226_ b_h\[11\] VGND VGND VPWR VPWR _09646_ sky130_fd_sc_hd__inv_16
XPHY_EDGE_ROW_144_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18871_ _09747_ _09760_ _09761_ VGND VGND VPWR VPWR _09763_ sky130_fd_sc_hd__nand3_1
X_17822_ _08679_ _08680_ _08675_ VGND VGND VPWR VPWR _08683_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17753_ _08543_ _08460_ _08457_ _08456_ VGND VGND VPWR VPWR _08616_ sky130_fd_sc_hd__nand4_1
X_14965_ _05819_ _05820_ _05857_ _05858_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a22o_1
X_16704_ net237 _07573_ _07574_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__nand3b_2
X_17684_ _08474_ _08476_ _08524_ VGND VGND VPWR VPWR _08547_ sky130_fd_sc_hd__o21ai_1
XFILLER_75_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13916_ _04680_ _04700_ _04816_ _04817_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__o211ai_2
X_16635_ _07506_ _07503_ _07492_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__a21o_1
X_14896_ net750 net642 VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__nand2_1
X_19423_ _00602_ _00598_ _00594_ _00603_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__o211a_1
XFILLER_90_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13847_ _04592_ _04595_ _04597_ _04753_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__o211ai_4
XFILLER_35_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16566_ _07060_ _07437_ _07436_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__a21o_1
X_13778_ _04585_ net211 VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__nand2_1
XFILLER_43_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19354_ _00530_ _00531_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__nand2_1
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16497_ _07241_ _07368_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__nand2_1
X_15517_ net627 net1105 _09581_ _09166_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__o2bb2a_1
X_18305_ _09150_ _09151_ VGND VGND VPWR VPWR _09152_ sky130_fd_sc_hd__nand2_1
X_12729_ _03630_ _03632_ _03655_ VGND VGND VPWR VPWR _03659_ sky130_fd_sc_hd__o21ai_1
X_19285_ _00455_ _00456_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__nand2_2
XFILLER_30_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18236_ _09077_ _09046_ _09076_ VGND VGND VPWR VPWR _09083_ sky130_fd_sc_hd__nand3_4
X_15448_ _06302_ _06338_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__nand2_1
X_18167_ _09011_ _09012_ _08895_ _08896_ VGND VGND VPWR VPWR _09015_ sky130_fd_sc_hd__o2bb2ai_1
X_15379_ _06229_ _06269_ _06270_ _06095_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__nand4b_2
Xhold426 p_hh\[16\] VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 p_hh\[24\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17118_ _07983_ _07984_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__nand2_4
X_18098_ _08831_ _08887_ _08940_ _08942_ _08885_ VGND VGND VPWR VPWR _08947_ sky130_fd_sc_hd__a221o_1
Xhold404 p_ll_pipe\[19\] VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold437 p_hh_pipe\[14\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap145 _07436_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_132_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold448 term_low\[2\] VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ _07912_ _07898_ _07916_ VGND VGND VPWR VPWR _07918_ sky130_fd_sc_hd__o21ai_1
Xhold459 p_ll\[16\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap189 _08951_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
X_20060_ _01288_ _01291_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__nand2_1
XFILLER_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_129_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_142_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20327_ net794 net25 VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__and2_1
XFILLER_135_699 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11060_ net678 net547 VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__nand2_1
XFILLER_1_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap690 a_h\[5\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__buf_6
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20258_ _09351_ _09373_ _01412_ _01463_ _01466_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__o311a_1
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20189_ _01358_ _01378_ _01379_ _01427_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14750_ _05643_ _05645_ _05549_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__a21o_1
X_11962_ _02738_ _02896_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__nand2_4
XFILLER_56_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13701_ _02082_ net922 VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__nor2_4
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11893_ _02828_ net475 net708 VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__and3_1
X_10913_ net707 net702 net441 _01861_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a31oi_1
X_14681_ net425 _05577_ _05566_ _05567_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__a211o_1
X_16420_ _07081_ _07085_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__nand2_1
X_10844_ net795 net1158 VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__and2_1
X_13632_ _04540_ _04530_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nand2_1
X_16351_ _07120_ _07107_ _07109_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__o21ai_1
X_13563_ _04396_ _04464_ _04470_ _04373_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__a211o_1
X_10775_ _01794_ _01798_ _01800_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__o21a_1
X_12514_ _03262_ _03441_ _03440_ net354 VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__o211a_1
X_19070_ _09924_ _09959_ VGND VGND VPWR VPWR _09961_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ _06194_ net224 net715 net944 VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__nand4_4
X_16282_ _07155_ _07156_ VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__nand2_2
X_18021_ net790 net605 VGND VGND VPWR VPWR _08871_ sky130_fd_sc_hd__nand2_1
X_13494_ net773 net766 net689 net683 VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__nand4_2
X_12445_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15233_ _06047_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__nor2_1
X_12376_ net679 net489 VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15164_ _06058_ _06060_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__nand2_1
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11327_ _02192_ _02197_ _02263_ _02264_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__a22o_1
X_14115_ net981 _05018_ _05009_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__and3_1
XFILLER_4_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19972_ _01193_ _01195_ _09253_ _09384_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__o2bb2ai_2
X_15095_ _05942_ _05947_ _05957_ _05990_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__o211ai_1
XFILLER_141_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11258_ _02196_ _02191_ _02188_ _02195_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__o211ai_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14046_ _04835_ _04948_ _04949_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__nand3_2
X_18923_ _09812_ _09813_ VGND VGND VPWR VPWR _09815_ sky130_fd_sc_hd__nand2_1
X_11189_ _02120_ _02121_ _02125_ _02043_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__a31oi_2
X_10209_ net867 VGND VGND VPWR VPWR _09460_ sky130_fd_sc_hd__inv_8
X_18854_ net630 net721 _09743_ _09744_ VGND VGND VPWR VPWR _09746_ sky130_fd_sc_hd__a22o_1
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17805_ _08664_ _08665_ _08666_ VGND VGND VPWR VPWR _08667_ sky130_fd_sc_hd__a21oi_1
X_15997_ _06873_ _06859_ _06872_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__nand3_4
X_18785_ _09637_ _09674_ _09673_ VGND VGND VPWR VPWR _09676_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_124_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17736_ _08596_ _08597_ net1072 net472 VGND VGND VPWR VPWR _08599_ sky130_fd_sc_hd__nand4_2
XFILLER_48_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14948_ _05679_ _05686_ _05687_ _05696_ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__a31oi_2
XFILLER_36_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17667_ _08443_ _08430_ _08429_ VGND VGND VPWR VPWR _08531_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14879_ _05658_ _05666_ _05778_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__a21oi_1
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16618_ _07367_ _07408_ _07405_ _07400_ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_106_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17598_ _08458_ _08462_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__nor2_1
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19406_ _00586_ _00587_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__nor2_2
X_16549_ _07348_ _07415_ _07416_ _07287_ _07285_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__a32oi_2
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19337_ net618 net718 _00509_ _00510_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_139_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19268_ net919 net552 VGND VGND VPWR VPWR _10170_ sky130_fd_sc_hd__nand2_2
X_18219_ net791 net782 net593 net585 VGND VGND VPWR VPWR _09066_ sky130_fd_sc_hd__nand4_4
X_19199_ _10089_ net732 net603 VGND VGND VPWR VPWR _10096_ sky130_fd_sc_hd__nand3_1
XFILLER_132_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20112_ _01179_ _01272_ _01269_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__o21a_1
X_20043_ _01270_ net143 _01269_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__o21ai_1
XFILLER_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10560_ net793 net1191 VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__and2_1
X_10491_ _01645_ term_high\[50\] term_high\[49\] net1367 VGND VGND VPWR VPWR _01649_
+ sky130_fd_sc_hd__a31o_1
XFILLER_139_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer320 net587 VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_147_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12230_ _03162_ _03163_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer353 net1149 VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12161_ net983 net474 _03094_ _03095_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__a22oi_2
XFILLER_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11112_ _02052_ _02053_ _01984_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__a21boi_4
X_12092_ _03025_ _03021_ _03024_ net1034 VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_92_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ _01979_ _01981_ _01984_ _01985_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__o2bb2ai_2
X_15920_ _06793_ _06794_ _06797_ _06658_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_104_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15851_ _06727_ net173 VGND VGND VPWR VPWR _06730_ sky130_fd_sc_hd__nand2_1
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14802_ _05698_ _05677_ _05697_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__nand3_2
X_15782_ net624 net628 net512 net505 VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__nand4_2
X_18570_ _09322_ _09441_ VGND VGND VPWR VPWR _09442_ sky130_fd_sc_hd__nand2_1
X_12994_ _03918_ _03728_ _03917_ VGND VGND VPWR VPWR _03921_ sky130_fd_sc_hd__nand3_1
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11945_ _02742_ _02743_ _02731_ _02729_ _02728_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a32oi_4
X_17521_ net1093 net485 net479 net581 VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__a22o_1
X_14733_ net285 _05599_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__nand2_1
XFILLER_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ net581 net485 net479 net585 VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__a22o_1
XFILLER_44_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14664_ _05418_ _05422_ _05421_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__a21bo_2
XFILLER_33_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11876_ _02688_ _02811_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__and2_1
X_16403_ _07270_ _07272_ _07259_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__a21oi_1
X_13615_ _04521_ _04522_ _04517_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__a21o_1
XFILLER_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17383_ _08247_ _08248_ VGND VGND VPWR VPWR _08250_ sky130_fd_sc_hd__nand2_1
X_10827_ p_hl\[29\] p_lh\[29\] _01844_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__a21o_1
X_14595_ net349 _05358_ _05494_ _05495_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_15_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16334_ _07199_ _07202_ _07205_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__a21o_1
X_10758_ _01759_ _01783_ _01782_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__a21oi_1
X_13546_ _04452_ _04453_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__nand2_2
X_19122_ _09939_ _09943_ _09940_ VGND VGND VPWR VPWR _10012_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16265_ _06901_ _06958_ _09188_ _09613_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_101_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13477_ net165 _04386_ _04387_ _09690_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__o211a_1
X_19053_ _09941_ _09943_ _09220_ _09286_ VGND VGND VPWR VPWR _09944_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12428_ _03225_ net474 net706 _03223_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__a31o_1
X_18004_ net338 net306 _08854_ VGND VGND VPWR VPWR _08855_ sky130_fd_sc_hd__a21o_1
X_10689_ p_hl\[9\] p_lh\[9\] _01726_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__o21a_1
X_15216_ _06110_ net669 net719 _06109_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__and4_1
X_16196_ net842 net620 net496 net491 _07066_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__a41o_1
XFILLER_138_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12359_ _03272_ _03274_ _03289_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o21ai_1
X_15147_ _06006_ _06037_ _06040_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__nand3_1
X_19955_ _01085_ _01173_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__nand2_1
X_15078_ net1055 _05865_ _05871_ _05972_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__o211ai_4
XFILLER_113_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14029_ _04933_ _04918_ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__nand2_1
X_18906_ net763 net580 VGND VGND VPWR VPWR _09798_ sky130_fd_sc_hd__nand2_1
X_19886_ _01101_ _01102_ VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__or2_1
X_18837_ _09729_ _09725_ VGND VGND VPWR VPWR _09730_ sky130_fd_sc_hd__nand2_1
XFILLER_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18768_ net792 net560 VGND VGND VPWR VPWR _09658_ sky130_fd_sc_hd__nand2_1
X_17719_ _08562_ _08575_ _08576_ _08377_ VGND VGND VPWR VPWR _08582_ sky130_fd_sc_hd__a31oi_1
X_20730_ clknet_leaf_36_clk _00370_ VGND VGND VPWR VPWR p_ll\[0\] sky130_fd_sc_hd__dfxtp_1
X_18699_ _09443_ _09576_ _09577_ VGND VGND VPWR VPWR _09583_ sky130_fd_sc_hd__nand3_1
XFILLER_51_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20661_ clknet_leaf_12_clk _00301_ VGND VGND VPWR VPWR p_hh\[27\] sky130_fd_sc_hd__dfxtp_1
X_20592_ clknet_leaf_12_clk _00232_ VGND VGND VPWR VPWR p_hh_pipe\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_750 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20026_ _01251_ _01252_ _01152_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__a21oi_1
XFILLER_86_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11730_ _02519_ _02540_ _02517_ _02520_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__o2bb2ai_2
Xrebuffer60 net856 VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__buf_2
Xrebuffer71 a_h\[12\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_15_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer82 net878 VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__buf_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer93 _03953_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__clkbuf_2
X_11661_ _02575_ _02594_ _02595_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__nand3b_1
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11592_ _02528_ _02529_ _02530_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__a21oi_1
X_13400_ _04310_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__nand2_1
X_10612_ net794 net1216 VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ net778 net639 VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__nand2_1
X_10543_ net793 net1234 VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__and2_1
X_13331_ _04242_ _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__nand2_1
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16050_ _06917_ _06923_ _06855_ _06922_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__o211ai_4
Xrebuffer150 net545 VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_77_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10474_ term_mid\[48\] term_high\[48\] VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__and2_1
Xrebuffer183 net654 VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlymetal6s2s_1
X_13262_ _04143_ _04154_ _04174_ _04175_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__a22o_1
X_15001_ _05838_ _05840_ _05853_ _05898_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__o211ai_2
Xrebuffer161 net957 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__buf_1
XFILLER_142_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer194 _02042_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12213_ _02738_ net535 net633 VGND VGND VPWR VPWR _03147_ sky130_fd_sc_hd__and3_1
X_13193_ _04087_ _04094_ _04112_ _04086_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__o211ai_1
X_12144_ _02831_ _02844_ _03068_ net268 _02843_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_90_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19740_ _00808_ _00813_ _00939_ _00940_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__a22o_1
X_12075_ net644 net526 net1059 net647 VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__a22oi_1
X_16952_ net566 net558 net523 net516 VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__and4_2
X_15903_ _06774_ _06775_ _06771_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__a21o_1
X_11026_ _01965_ _01966_ _01957_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__a21oi_1
X_16883_ _07750_ _07751_ VGND VGND VPWR VPWR _07753_ sky130_fd_sc_hd__nand2_1
X_19671_ net877 net553 VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__nand2_1
X_15834_ _06709_ _06710_ _06672_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__and3_1
X_18622_ net763 net596 VGND VGND VPWR VPWR _09498_ sky130_fd_sc_hd__nand2_1
XFILLER_49_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18553_ _09402_ _09403_ _09421_ VGND VGND VPWR VPWR _09423_ sky130_fd_sc_hd__a21oi_1
X_15765_ _06643_ _06644_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__nand2_1
X_17504_ _08270_ _08282_ _08368_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__and3_1
X_12977_ net1049 net824 VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__nand2_2
X_15696_ _06511_ _06553_ _06554_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__a21oi_1
X_11928_ net665 net508 VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__nand2_1
X_18484_ _09270_ _09273_ _09276_ _09343_ _09344_ VGND VGND VPWR VPWR _09347_ sky130_fd_sc_hd__o2111a_1
X_14716_ net740 net736 net670 net668 VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__nand4_1
X_11859_ _02793_ _02794_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__nand2_1
X_17435_ _08176_ _08188_ _08178_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__o21a_2
X_14647_ _05544_ _05545_ net716 net699 VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_31_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_29 net487 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _00436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17366_ net234 _08232_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__nand2_1
X_14578_ _05347_ _05479_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__nand2_1
X_16317_ net620 net491 VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_119_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19105_ _09991_ _09995_ _09736_ VGND VGND VPWR VPWR _09996_ sky130_fd_sc_hd__a21o_1
X_13529_ net748 net711 VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nand2_1
X_17297_ _07992_ _08134_ _08137_ _08139_ _08040_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__a32oi_2
X_16248_ _07108_ _07109_ _07120_ VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__and3_1
X_19036_ _09811_ _09817_ _09814_ VGND VGND VPWR VPWR _09927_ sky130_fd_sc_hd__a21o_1
Xoutput103 net103 VGND VGND VPWR VPWR p[43] sky130_fd_sc_hd__buf_2
Xoutput114 net114 VGND VGND VPWR VPWR p[53] sky130_fd_sc_hd__buf_2
Xoutput125 net125 VGND VGND VPWR VPWR p[63] sky130_fd_sc_hd__buf_2
X_16179_ _06841_ _06941_ _06948_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_132_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19938_ _01094_ _01096_ _01157_ _01158_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__nand4_2
XFILLER_68_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19869_ _01055_ _01065_ _01054_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_147_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20713_ clknet_leaf_55_clk net132 VGND VGND VPWR VPWR p_lh\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_12_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20644_ clknet_leaf_17_clk _00284_ VGND VGND VPWR VPWR p_hh\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20575_ clknet_leaf_27_clk _00215_ VGND VGND VPWR VPWR p_hh_pipe\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10190_ net588 VGND VGND VPWR VPWR _09253_ sky130_fd_sc_hd__inv_8
XFILLER_2_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_127_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone109 net980 VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__clkbuf_16
XFILLER_59_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12900_ net645 net638 net856 net823 VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__nand4_1
X_13880_ _04661_ _04664_ _04662_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__a21oi_1
X_20009_ _01232_ _01233_ _01215_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__a21oi_2
X_12831_ net396 _03754_ _03756_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_87_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15550_ net631 net611 net1041 net522 VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__and4_1
X_12762_ _03620_ _03622_ _03690_ _03691_ VGND VGND VPWR VPWR _03692_ sky130_fd_sc_hd__o211ai_1
X_11713_ net682 net679 net511 net508 VGND VGND VPWR VPWR _02651_ sky130_fd_sc_hd__nand4_2
X_12693_ net682 net474 _03618_ _03619_ VGND VGND VPWR VPWR _03623_ sky130_fd_sc_hd__a22o_1
XFILLER_14_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14501_ _05111_ _05113_ _05399_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__o21a_1
X_15481_ net716 _06264_ _06370_ net722 VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__o22a_1
X_11644_ _02579_ _02580_ _02578_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__o21bai_1
X_17220_ _07971_ _07972_ _07964_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__o21ai_1
X_14432_ net720 net703 VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__and2_1
X_17151_ _08012_ _08014_ _08019_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__a21o_1
XFILLER_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput27 a[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
X_16102_ _06861_ _06864_ _06869_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__o21ai_1
X_11575_ _02483_ _02489_ _02490_ net359 _02512_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__o2111ai_4
X_14363_ _05119_ _05238_ _05240_ _05245_ _05116_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__a32oi_4
Xwire742 b_l\[9\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__buf_12
Xinput16 a[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_10526_ term_high\[61\] term_high\[62\] _01669_ net1310 VGND VGND VPWR VPWR _01672_
+ sky130_fd_sc_hd__a31oi_1
X_17082_ net593 net488 VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__and2_1
Xmax_cap508 net509 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__buf_12
X_13314_ _04225_ net693 net777 _04223_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__nand4_1
Xinput49 b[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 b[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
X_14294_ _05194_ _05196_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__nor2_1
Xwire764 net765 VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__buf_6
X_10457_ term_mid\[44\] term_high\[44\] _01619_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__a21bo_1
X_16033_ net624 net1045 net512 net505 _06791_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__a41o_1
XFILLER_109_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap519 net520 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__buf_12
X_13245_ _04148_ net710 net777 _04146_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__a31o_1
XFILLER_6_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10388_ term_mid\[35\] term_high\[35\] VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__xor2_1
X_13176_ net641 b_h\[15\] VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__nand2_1
X_12127_ _03059_ net461 _03049_ _03058_ VGND VGND VPWR VPWR _03062_ sky130_fd_sc_hd__o211ai_4
XFILLER_111_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17984_ _08819_ net779 net628 _08820_ VGND VGND VPWR VPWR _08835_ sky130_fd_sc_hd__a31oi_1
X_12058_ _02986_ _02989_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__nand2_1
X_16935_ _07802_ _07804_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__nand2_1
XFILLER_78_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19723_ _00929_ _00923_ _00928_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__and3_1
X_11009_ _01952_ _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nand2_1
XFILLER_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19654_ _00708_ _00716_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__nand2_1
X_16866_ _07678_ _07683_ _07679_ _07674_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__o2bb2ai_2
X_18605_ net792 net564 VGND VGND VPWR VPWR _09479_ sky130_fd_sc_hd__nand2_1
XFILLER_53_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15817_ _06693_ _06694_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__nand2_2
X_16797_ net572 net513 VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__nand2_1
XFILLER_18_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19585_ _00459_ _00663_ _00661_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__o21ai_1
X_15748_ net383 _06583_ _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__o21ai_1
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18536_ net621 net743 VGND VGND VPWR VPWR _09404_ sky130_fd_sc_hd__nand2_1
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18467_ _09248_ _09249_ _09251_ VGND VGND VPWR VPWR _09328_ sky130_fd_sc_hd__o21a_1
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15679_ _06554_ _06556_ _06557_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__o21ai_1
X_17418_ _08243_ _08241_ _08240_ _08259_ VGND VGND VPWR VPWR _08284_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_44_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18398_ net604 net764 _09250_ _09251_ VGND VGND VPWR VPWR _09254_ sky130_fd_sc_hd__a22o_1
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17349_ _09319_ _09613_ _08211_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__o21ai_1
X_20360_ clknet_leaf_51_clk _00000_ VGND VGND VPWR VPWR b_l\[0\] sky130_fd_sc_hd__dfxtp_4
X_20291_ _01505_ _01506_ _01532_ _01533_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__nor4_1
X_19019_ _09908_ _09909_ VGND VGND VPWR VPWR _09910_ sky130_fd_sc_hd__nand2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20627_ clknet_leaf_47_clk _00267_ VGND VGND VPWR VPWR p_ll_pipe\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20558_ clknet_leaf_27_clk _00198_ VGND VGND VPWR VPWR mid_sum\[21\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11360_ _02295_ _02299_ _02297_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a21oi_1
XFILLER_118_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10311_ _00784_ _00795_ _00773_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__a21oi_1
X_20489_ clknet_leaf_28_clk _00129_ VGND VGND VPWR VPWR term_mid\[33\] sky130_fd_sc_hd__dfxtp_1
X_11291_ net201 _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__nand2_1
XFILLER_98_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13030_ net793 _03955_ _03956_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__and3_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10242_ net794 net35 VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__and2_1
XFILLER_79_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_120_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16720_ _07489_ _07557_ _07554_ _07550_ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_89_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14981_ _05755_ _05758_ _05873_ _05874_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a22o_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13932_ net724 net709 net431 _04836_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a31oi_2
X_16651_ net876 net541 VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__and2_1
XFILLER_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13863_ _04723_ _04726_ _04767_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__o21ai_2
XFILLER_19_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16582_ _07352_ _07362_ _07364_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__o21a_1
X_15602_ net1070 _06480_ net612 net540 _06479_ VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__o2111ai_4
XFILLER_90_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12814_ _09635_ _03639_ _03636_ _03641_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__o22a_1
X_13794_ _04563_ _04681_ _04684_ _04686_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__o2bb2ai_4
X_19370_ _00546_ net230 _00545_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__a21oi_1
X_15533_ _09144_ _09581_ _06414_ _06416_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__o211a_1
X_18321_ _09164_ _09160_ _09133_ _09165_ VGND VGND VPWR VPWR _09170_ sky130_fd_sc_hd__o211ai_4
X_12745_ _03672_ _03673_ net645 b_h\[8\] VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__nand4_1
XFILLER_42_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12676_ _03373_ _03371_ _03495_ _03247_ _03606_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a41oi_2
X_18252_ net187 net207 _09094_ VGND VGND VPWR VPWR _09099_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_41_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _06347_ _06348_ _06353_ _06354_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__nor4_1
X_11627_ _02564_ _02560_ _02563_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__a21o_1
X_17203_ _08060_ _08065_ _08069_ _08063_ VGND VGND VPWR VPWR _08071_ sky130_fd_sc_hd__o211ai_1
X_18183_ _09029_ net749 net630 _09028_ VGND VGND VPWR VPWR _09030_ sky130_fd_sc_hd__nand4_4
X_15395_ _06283_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__nor2_1
X_14415_ _05312_ _05313_ _05314_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_116_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17134_ _07896_ _07997_ _07895_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__a21oi_2
X_11558_ net658 net535 VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__nand2_1
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14346_ _05116_ _05242_ _05245_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__nand3b_4
XFILLER_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10509_ net1356 _01660_ _01661_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__o21a_1
Xwire583 net584 VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__buf_12
X_17065_ _07930_ _07822_ _07929_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__nand3_2
Xmax_cap305 _08898_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_1
X_11489_ _02423_ _02424_ net269 VGND VGND VPWR VPWR _02429_ sky130_fd_sc_hd__a21o_1
X_16016_ _06768_ _06856_ _06891_ _06892_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__o211a_1
Xmax_cap338 _08818_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlymetal6s2s_1
Xmax_cap349 _05353_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_2
X_14277_ _05143_ _05178_ _05176_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13228_ net713 net923 VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__nand2_1
XFILLER_124_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13159_ _04081_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__inv_2
X_17967_ net623 net781 net615 net790 VGND VGND VPWR VPWR _08819_ sky130_fd_sc_hd__a22o_1
X_19706_ net580 b_l\[11\] VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_144_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16918_ _07783_ _07786_ _09275_ _09613_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__o2bb2ai_1
X_17898_ _08755_ _08756_ VGND VGND VPWR VPWR _08757_ sky130_fd_sc_hd__nand2_1
X_16849_ _07715_ _07717_ _07588_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__nand3_1
XFILLER_81_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19637_ _00829_ _00834_ _00836_ _00729_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__o211ai_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19568_ _09264_ _09286_ _00651_ _00653_ _00455_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__o32a_1
X_18519_ _09385_ _09353_ _09383_ VGND VGND VPWR VPWR _09386_ sky130_fd_sc_hd__nand3_4
XFILLER_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19499_ _10160_ _00486_ _00528_ _00529_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__a22oi_1
X_20412_ clknet_leaf_30_clk _00052_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20343_ net793 net7 VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__and2_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20274_ _01437_ _01477_ _01479_ _01480_ _01483_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__a32oi_2
XTAP_TAPCELL_ROW_8_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10860_ net793 net1260 VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__and2_1
XFILLER_56_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10791_ _01808_ _01814_ net796 VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__a21oi_1
X_12530_ _03295_ _03378_ _03458_ _03459_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__a22oi_1
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12461_ _09624_ _03388_ net489 net674 _03387_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__o2111ai_4
XFILLER_138_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11412_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__inv_2
X_14200_ _05098_ _05103_ _05100_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__or3b_4
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15180_ _06070_ _06072_ _06075_ _05890_ _06074_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__a221oi_1
XFILLER_126_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12392_ _03304_ _03305_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__o21ai_1
X_14131_ _05004_ _05006_ _05026_ _05028_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__o2bb2ai_1
X_11343_ _09460_ _09592_ _01857_ _02278_ _02277_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__o221ai_4
X_11274_ _02215_ _02214_ _02150_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_111_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14062_ _04869_ _04945_ _04940_ _04946_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__o2bb2ai_1
X_10225_ net495 VGND VGND VPWR VPWR _09635_ sky130_fd_sc_hd__inv_6
X_13013_ _03938_ _03939_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__nand2_1
X_18870_ _09760_ _09761_ _09747_ VGND VGND VPWR VPWR _09762_ sky130_fd_sc_hd__a21o_1
X_17821_ _08629_ _08676_ a_l\[12\] net477 _08680_ VGND VGND VPWR VPWR _08682_ sky130_fd_sc_hd__o2111ai_4
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17752_ _08456_ _08457_ _08541_ _08542_ VGND VGND VPWR VPWR _08615_ sky130_fd_sc_hd__nand4_4
XFILLER_66_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14964_ _05819_ _05820_ _05857_ _05858_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nand4_1
X_16703_ _07573_ _07574_ net237 VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__a21bo_1
X_17683_ _08545_ _08463_ net795 _08546_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__o211a_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13915_ _04700_ _04680_ _04816_ net164 VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__o211a_4
X_16634_ net453 _07394_ _07504_ _07505_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__o211ai_4
XFILLER_90_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19422_ _00599_ _00601_ _00595_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__a21o_1
X_14895_ net756 net1135 VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__nand2_1
X_13846_ _02502_ _04134_ _04743_ _04747_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__o211ai_2
X_16565_ _07437_ _07060_ VGND VGND VPWR VPWR _07438_ sky130_fd_sc_hd__nand2_4
X_10989_ _01933_ _01934_ _01883_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__a21boi_1
X_13777_ _04655_ _04660_ _04675_ _04676_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_31_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19353_ _00524_ _00525_ _00527_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__nand3_1
X_16496_ _07227_ _07236_ _07237_ _07251_ _07240_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__a32oi_2
X_15516_ net627 net631 VGND VGND VPWR VPWR _06402_ sky130_fd_sc_hd__nand2_8
X_18304_ net791 net782 net585 net582 VGND VGND VPWR VPWR _09151_ sky130_fd_sc_hd__nand4_4
X_12728_ _03631_ _03633_ _03652_ _03653_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__nand4_1
X_19284_ net754 net575 net567 net760 VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__a22oi_1
X_12659_ _03574_ _03575_ _03503_ _03585_ _03586_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__a32oi_4
X_18235_ _09047_ _09078_ _09079_ VGND VGND VPWR VPWR _09082_ sky130_fd_sc_hd__nand3_4
X_15447_ _06301_ _06334_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__and2b_1
XFILLER_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_128_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18166_ _09011_ _09012_ _08898_ VGND VGND VPWR VPWR _09014_ sky130_fd_sc_hd__nand3_1
X_15378_ net730 _06095_ net635 _06270_ _06269_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__a32o_1
Xwire380 _07032_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold427 mid_sum\[18\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 p_hh_pipe\[1\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
X_17117_ _07761_ _07768_ _07978_ _07982_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__o211ai_2
X_18097_ _08940_ _08942_ _08944_ VGND VGND VPWR VPWR _08946_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold416 p_ll_pipe\[22\] VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ _05223_ _05224_ _05226_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__a21o_1
Xwire391 _05164_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_1
Xhold438 p_hh_pipe\[11\] VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap146 net147 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
X_17048_ _07898_ _07912_ _07916_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__o21a_1
Xhold449 p_ll_pipe\[20\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap168 _01538_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18999_ _09884_ net852 _09880_ _09888_ VGND VGND VPWR VPWR _09890_ sky130_fd_sc_hd__o211ai_4
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone281 net687 VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__clkbuf_16
XFILLER_93_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20326_ net794 net24 VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__and2_1
XFILLER_134_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap691 net692 VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__buf_12
XFILLER_1_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap680 a_h\[7\] VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__buf_12
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20257_ _01498_ _01350_ _01501_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__a21oi_4
XFILLER_135_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20188_ _01358_ _01378_ _01379_ _01427_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__a31oi_2
XFILLER_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11961_ net633 net546 net537 net1036 VGND VGND VPWR VPWR _02897_ sky130_fd_sc_hd__a22oi_4
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10912_ net702 net947 net538 net707 VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__a22oi_1
XFILLER_57_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13700_ net768 net676 net673 net773 VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__a22oi_4
X_11892_ net706 net698 net483 net481 VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__nand4_1
XFILLER_45_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14680_ _05568_ _05578_ _05579_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__nand3_1
X_10843_ net795 net1190 VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__and2_1
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13631_ _04513_ _04515_ _04533_ _04531_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__a22oi_2
X_16350_ _07149_ net280 _07126_ _07123_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__o2bb2ai_1
X_10774_ _01792_ _01793_ _01797_ net795 VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__o31a_1
X_13562_ _04470_ _04373_ _04469_ _04468_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__o211ai_2
X_16281_ _07152_ _07089_ _07153_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__nand3_4
X_12513_ _03439_ _03440_ _03442_ _03259_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15301_ _06194_ net224 _09384_ _09471_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__o2bb2ai_2
X_18020_ net781 net886 VGND VGND VPWR VPWR _08870_ sky130_fd_sc_hd__nand2_1
X_13493_ net773 net683 VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__nand2_1
XFILLER_12_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12444_ _03350_ _03353_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15232_ _06126_ _06127_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__nand2_1
XFILLER_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12375_ _03187_ _03188_ _03185_ VGND VGND VPWR VPWR _03308_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_10_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15163_ _06055_ _06049_ _05989_ _06057_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__o211ai_2
XFILLER_126_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11326_ _02263_ _02264_ _02265_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__a21bo_1
XFILLER_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19971_ _09253_ _09384_ _01193_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__o21ai_1
X_15094_ _05942_ _05947_ _05957_ _05990_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__o211a_1
X_14114_ _04876_ net430 _05015_ _05016_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__o211ai_4
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18922_ net817 net557 net1102 net1057 VGND VGND VPWR VPWR _09814_ sky130_fd_sc_hd__a22oi_4
X_14045_ _04862_ _04867_ _04868_ _04945_ _04947_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__o2111ai_4
X_11257_ _02191_ _02197_ _02187_ _02198_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__o211ai_4
XFILLER_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11188_ _02126_ _02128_ _02040_ _02041_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__o2bb2ai_2
X_10208_ net680 VGND VGND VPWR VPWR _09449_ sky130_fd_sc_hd__inv_8
X_18853_ _05044_ _06441_ net630 net721 _09743_ VGND VGND VPWR VPWR _09745_ sky130_fd_sc_hd__o2111ai_2
Xsplit122 b_l\[4\] VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__clkbuf_4
XFILLER_121_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17804_ _08607_ _08610_ VGND VGND VPWR VPWR _08666_ sky130_fd_sc_hd__nand2_1
X_18784_ _09671_ _09672_ VGND VGND VPWR VPWR _09675_ sky130_fd_sc_hd__nand2_1
X_15996_ _06864_ _06868_ _06861_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__o21ai_1
X_17735_ net1072 net472 _08596_ _08597_ VGND VGND VPWR VPWR _08598_ sky130_fd_sc_hd__a22o_1
XFILLER_36_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14947_ _05844_ _05834_ _05833_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__nand3_1
XFILLER_36_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17666_ _08475_ _08477_ _08524_ _08526_ VGND VGND VPWR VPWR _08530_ sky130_fd_sc_hd__nand4_1
XFILLER_63_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14878_ _05775_ _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__nand2_1
X_16617_ _07486_ _07488_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_106_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17597_ _08280_ _08461_ _08460_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__a21oi_2
X_13829_ net762 net676 _04732_ _04734_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__a22oi_4
X_19405_ _00585_ _00580_ _00583_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__and3_4
X_16548_ _07417_ net208 _07310_ _07418_ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_18_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19336_ net618 net718 _00509_ _00510_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_139_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16479_ _07129_ _07262_ _07267_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__o21a_1
X_19267_ net808 net556 net552 net776 VGND VGND VPWR VPWR _10168_ sky130_fd_sc_hd__a22o_1
X_18218_ net791 net782 net593 net585 VGND VGND VPWR VPWR _09065_ sky130_fd_sc_hd__and4_1
X_19198_ _09885_ net927 _10090_ _10093_ VGND VGND VPWR VPWR _10095_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_129_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18149_ _08980_ _08982_ _08989_ _08991_ VGND VGND VPWR VPWR _08997_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_116_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20111_ _01182_ _01183_ _01273_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nand3_2
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20042_ _01270_ net143 _01269_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__o21a_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10490_ _01647_ _01648_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__nor2_1
Xrebuffer310 _06908_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__buf_2
Xrebuffer321 _09012_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlymetal6s4s_1
Xrebuffer332 _04544_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__clkbuf_2
XFILLER_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer354 net1149 VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlymetal6s2s_1
X_12160_ _03091_ _02856_ _02851_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__nand3b_1
X_11111_ _01982_ _01983_ _02052_ _02053_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__o211a_4
XFILLER_122_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12091_ _02906_ _02909_ _03019_ _03020_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__nand4_1
X_20309_ _01553_ _01550_ net794 _01555_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__o211a_1
XFILLER_1_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ _01980_ _01975_ net1075 _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__o211ai_2
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15850_ net191 _06652_ _06722_ _06723_ VGND VGND VPWR VPWR _06729_ sky130_fd_sc_hd__o211ai_2
XFILLER_103_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14801_ _05698_ _05677_ _05697_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__and3_1
X_15781_ net624 net628 net512 net505 VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__and4_1
X_12993_ _03896_ _03898_ _03914_ _03916_ VGND VGND VPWR VPWR _03920_ sky130_fd_sc_hd__o211ai_1
XFILLER_18_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11944_ net324 _02878_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nor2_2
X_17520_ net581 net479 VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__nand2_1
X_14732_ _05600_ _05627_ _05628_ _05599_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__a31o_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11875_ _02688_ net146 VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__nor2_2
X_17451_ net448 _08314_ _08302_ _08315_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__o211ai_4
X_14663_ _05561_ net312 VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__nand2_1
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16402_ _07270_ _07272_ _07258_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__a21o_1
X_10826_ p_hl\[29\] p_lh\[29\] p_hl\[28\] p_lh\[28\] VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__o211a_1
X_13614_ _04521_ _04522_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__nand2_1
X_17382_ _08248_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__inv_2
XFILLER_60_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19121_ _09939_ _09943_ _09940_ VGND VGND VPWR VPWR _10011_ sky130_fd_sc_hd__a21o_1
X_14594_ net349 _05358_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_15_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16333_ _07199_ _07202_ net420 VGND VGND VPWR VPWR _07207_ sky130_fd_sc_hd__nand3_1
X_10757_ _01759_ _01783_ _01782_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__a21o_1
X_13545_ _04321_ _04324_ net352 _04451_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__and4_1
X_16264_ _06998_ _07004_ _07133_ _07136_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_101_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13476_ _04384_ _04318_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__nand2_2
X_10688_ _09559_ _09570_ _01716_ _01719_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__o211ai_2
X_19052_ net776 net810 net568 net564 VGND VGND VPWR VPWR _09943_ sky130_fd_sc_hd__nand4_2
X_12427_ _03359_ _03252_ _03358_ VGND VGND VPWR VPWR _03360_ sky130_fd_sc_hd__nand3_2
X_18003_ _08851_ _08853_ VGND VGND VPWR VPWR _08854_ sky130_fd_sc_hd__and2b_1
XFILLER_65_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15215_ net719 net944 _06109_ _06110_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__a22oi_2
X_16195_ _07067_ _07069_ _07066_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__o21ai_1
XFILLER_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12358_ _03273_ _03275_ _03287_ _03288_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__nand4_2
X_15146_ _06037_ _06040_ _06005_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__a21o_1
X_11309_ _02153_ _02182_ _02183_ _02213_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__a31oi_2
X_12289_ _03068_ _03078_ _03221_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__a21oi_1
X_19954_ _01085_ _01177_ _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__nand3b_4
X_15077_ _05894_ _05973_ _05974_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__nand3_2
XFILLER_141_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18905_ _09651_ _09667_ _09669_ VGND VGND VPWR VPWR _09797_ sky130_fd_sc_hd__a21boi_2
X_19885_ _01101_ _01102_ VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__nor2_1
X_14028_ _04933_ _04918_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__and2_1
XFILLER_110_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18836_ _09726_ _09722_ _09583_ VGND VGND VPWR VPWR _09729_ sky130_fd_sc_hd__a21oi_1
XFILLER_68_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15979_ _06766_ _06754_ _06765_ _06779_ _06781_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__a32oi_4
XFILLER_67_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18767_ net780 net568 VGND VGND VPWR VPWR _09656_ sky130_fd_sc_hd__nand2_1
X_17718_ _08575_ _08576_ _08562_ VGND VGND VPWR VPWR _08581_ sky130_fd_sc_hd__a21o_1
X_18698_ _09430_ _09433_ _09578_ _09579_ VGND VGND VPWR VPWR _09582_ sky130_fd_sc_hd__a22oi_1
XFILLER_36_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17649_ _08511_ _08512_ VGND VGND VPWR VPWR _08513_ sky130_fd_sc_hd__nand2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20660_ clknet_leaf_2_clk _00300_ VGND VGND VPWR VPWR p_hh\[26\] sky130_fd_sc_hd__dfxtp_1
X_20591_ clknet_leaf_12_clk _00231_ VGND VGND VPWR VPWR p_hh_pipe\[21\] sky130_fd_sc_hd__dfxtp_1
X_19319_ _10086_ _10089_ _10090_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__a21o_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20025_ _01152_ _01251_ net1029 VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__nand3_4
XFILLER_101_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer50 _06401_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_771 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer72 a_h\[12\] VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer61 net857 VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer94 a_h\[11\] VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer83 b_l\[6\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd1_1
X_11660_ _02596_ _02597_ _02575_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__a21oi_1
XFILLER_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11591_ _02373_ _02377_ _02375_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__a21oi_4
X_20789_ clknet_leaf_7_clk _00429_ VGND VGND VPWR VPWR a_l\[11\] sky130_fd_sc_hd__dfxtp_4
X_10611_ net794 net1254 VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ net793 net1204 VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__and2_1
XFILLER_128_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13330_ _04231_ _04232_ _04239_ _04240_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__nand4_2
Xrebuffer140 net936 VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd1_1
X_13261_ _04174_ _04175_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__nand2_1
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10473_ term_mid\[48\] term_high\[48\] VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__nor2_1
XFILLER_108_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer173 _07528_ VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__buf_2
Xrebuffer151 net947 VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlymetal6s2s_1
X_12212_ _03144_ _03145_ VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__nand2_1
X_15000_ _05850_ _05855_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__nand2_1
Xrebuffer162 net956 VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_136_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer195 _02042_ VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13192_ _04087_ _04094_ _04086_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__o21ai_1
Xrebuffer184 _05017_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__buf_4
X_12143_ _03069_ _03072_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__nand2_1
XFILLER_123_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16951_ net558 net516 VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__nand2_1
X_12074_ net647 net644 net526 net524 VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__nand4_2
X_15902_ _06774_ _06775_ _06771_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__a21oi_1
X_11025_ _01964_ _01969_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__nor2_2
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16882_ net586 net498 net493 net594 VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a22oi_2
XFILLER_77_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19670_ net819 net556 VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__nand2_1
X_15833_ _06710_ _06672_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__nand2_1
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18621_ net763 net596 VGND VGND VPWR VPWR _09497_ sky130_fd_sc_hd__and2_1
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15764_ _06640_ _06641_ _06564_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__nand3_4
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18552_ _09419_ _09420_ VGND VGND VPWR VPWR _09422_ sky130_fd_sc_hd__nor2_1
X_17503_ _08270_ _08282_ _08368_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__a21oi_1
X_12976_ net641 net826 VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__and2_1
X_14715_ net736 net668 VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__nand2_2
XFILLER_17_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15695_ _06555_ _06556_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _02707_ _02862_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__nand2_1
X_18483_ _09343_ _09344_ _09345_ VGND VGND VPWR VPWR _09346_ sky130_fd_sc_hd__a21boi_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11858_ _02793_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__and2_1
X_17434_ _08227_ _08296_ _08299_ VGND VGND VPWR VPWR _08300_ sky130_fd_sc_hd__o21a_1
X_14646_ _05544_ _05545_ _05541_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__and3_1
XFILLER_33_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10809_ _01827_ _01828_ _01829_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__o21a_1
X_11789_ net658 net653 net526 net520 VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__nand4_2
X_17365_ _08203_ _08226_ _08228_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__nand3_2
XANTENNA_19 _00437_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14577_ net740 net670 VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__nand2_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16316_ net841 net487 VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13528_ _01860_ _04260_ _04324_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__o21ai_2
X_19104_ _09867_ _09992_ _09993_ VGND VGND VPWR VPWR _09995_ sky130_fd_sc_hd__nand3_1
X_17296_ _08140_ _08146_ _08149_ _08144_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__o22ai_2
X_19035_ _09826_ _09831_ VGND VGND VPWR VPWR _09926_ sky130_fd_sc_hd__nand2_1
X_16247_ _07108_ _07109_ _07119_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__a21o_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13459_ _04333_ _04365_ _04366_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__nand3_1
Xoutput104 net104 VGND VGND VPWR VPWR p[44] sky130_fd_sc_hd__buf_2
Xoutput115 net115 VGND VGND VPWR VPWR p[54] sky130_fd_sc_hd__buf_2
X_16178_ _06833_ _06941_ _07052_ _07053_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__a31o_1
Xoutput126 net126 VGND VGND VPWR VPWR p[6] sky130_fd_sc_hd__buf_2
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15129_ _06021_ _06023_ _06018_ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__a21oi_1
XFILLER_101_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19937_ _01094_ _01096_ _01157_ _01158_ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a22o_1
XFILLER_96_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19868_ _01073_ _01068_ _01071_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_147_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18819_ _09630_ _09631_ _09707_ _09708_ VGND VGND VPWR VPWR _09712_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_39_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19799_ _01009_ _01011_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__nor2_1
XFILLER_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20712_ clknet_leaf_40_clk _00352_ VGND VGND VPWR VPWR p_lh\[14\] sky130_fd_sc_hd__dfxtp_1
X_20643_ clknet_leaf_17_clk _00283_ VGND VGND VPWR VPWR p_hh\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20574_ clknet_leaf_27_clk _00214_ VGND VGND VPWR VPWR p_hh_pipe\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20008_ _01215_ _01232_ _01233_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__nand3_2
XFILLER_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12830_ _03757_ _03741_ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__nand2_1
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12761_ _03681_ _03684_ _03685_ _03689_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__o211ai_4
XFILLER_55_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11712_ net679 net511 VGND VGND VPWR VPWR _02650_ sky130_fd_sc_hd__nand2_2
X_12692_ _03618_ _03619_ _03614_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__a21oi_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14500_ _05111_ _05113_ _05394_ _05399_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__a2bb2oi_4
X_15480_ net716 net640 VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__nand2_1
X_11643_ _01888_ _02338_ _02578_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__o21ai_1
X_14431_ net727 net1094 net699 net695 VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__nand4_4
X_17150_ _07868_ _07886_ _08018_ VGND VGND VPWR VPWR _08019_ sky130_fd_sc_hd__nand3_2
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 a[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
X_16101_ _06874_ _06975_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__nand2_1
X_11574_ net359 _02512_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__nand2_1
X_14362_ _05112_ b_l\[15\] net714 VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__and3_1
Xinput17 a[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
X_10525_ net1355 net1323 _01669_ _01671_ net65 VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__a311oi_1
X_17081_ _02338_ _06867_ _07749_ _07752_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__o22a_1
X_13313_ _04223_ _04225_ _09155_ _09417_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__o2bb2ai_1
Xmax_cap509 b_h\[7\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_12
Xinput39 b[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14293_ b_l\[14\] net709 _05192_ _05193_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__a22o_1
X_10456_ term_mid\[45\] term_high\[45\] VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__xor2_2
XFILLER_136_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16032_ net628 net502 _06658_ _06797_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__o2bb2a_1
X_13244_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__or2_1
XFILLER_6_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13175_ net634 b_h\[14\] VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__nand2_1
X_10387_ _01554_ _01559_ _01561_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__o21a_1
XFILLER_124_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12126_ net461 _03056_ _03048_ _03057_ VGND VGND VPWR VPWR _03061_ sky130_fd_sc_hd__o211ai_4
XFILLER_97_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17983_ net774 net769 _06401_ _08832_ VGND VGND VPWR VPWR _08834_ sky130_fd_sc_hd__a31o_1
XFILLER_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12057_ _02865_ _02866_ _02986_ _02988_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__a22o_1
X_16934_ net376 _07795_ _07799_ _07790_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__o211ai_1
X_19722_ _00920_ _00911_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__nand2_1
XFILLER_28_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11008_ _01949_ net517 net707 _01947_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__nand4_1
X_16865_ _07628_ _07695_ _07697_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__o21ai_1
X_19653_ _00853_ _00854_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__nand2_1
XFILLER_38_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15816_ net1117 net1041 net521 net613 VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__a22oi_1
XFILLER_92_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18604_ net782 net569 VGND VGND VPWR VPWR _09478_ sky130_fd_sc_hd__nand2_1
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16796_ net590 net503 VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__nand2_1
XFILLER_53_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19584_ _00777_ _00779_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__nand2_1
X_15747_ _06624_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__nand2_2
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12959_ _03881_ _03882_ _03879_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a21oi_1
X_18535_ _09399_ _09400_ _09325_ VGND VGND VPWR VPWR _09403_ sky130_fd_sc_hd__nand3_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15678_ _06553_ _06555_ _06510_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__a21o_1
X_18466_ _09248_ _09249_ _09251_ VGND VGND VPWR VPWR _09327_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17417_ _08243_ _08241_ _08240_ _08259_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__a22o_1
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14629_ _05395_ _05404_ _05527_ _05529_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__o22a_1
XFILLER_147_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18397_ _09250_ _09251_ _09210_ _09220_ VGND VGND VPWR VPWR _09252_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17348_ _08052_ _08210_ _08206_ _08208_ VGND VGND VPWR VPWR _08215_ sky130_fd_sc_hd__o211ai_2
X_17279_ net160 _08003_ _08141_ _08143_ VGND VGND VPWR VPWR _08147_ sky130_fd_sc_hd__o211ai_1
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20290_ _01505_ _01506_ _01532_ _01533_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__o22a_1
X_19018_ net758 net580 VGND VGND VPWR VPWR _09909_ sky130_fd_sc_hd__nand2_1
XFILLER_114_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20626_ clknet_leaf_48_clk _00266_ VGND VGND VPWR VPWR p_ll_pipe\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20557_ clknet_leaf_27_clk _00197_ VGND VGND VPWR VPWR mid_sum\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11290_ _02229_ _02149_ _02228_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__nand3_2
XFILLER_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10310_ term_low\[23\] term_mid\[23\] VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__or2_1
X_20488_ clknet_leaf_28_clk _00128_ VGND VGND VPWR VPWR term_mid\[32\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10241_ net794 net34 VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__and2_1
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14980_ _05755_ _05758_ _05873_ _05874_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_89_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13931_ _09177_ _09329_ _09351_ net709 VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__or4b_2
XFILLER_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16650_ _07372_ _07378_ _07375_ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__a21oi_2
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13862_ _04766_ _04767_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__nand2_1
XFILLER_35_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16581_ _07352_ _07362_ _07364_ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__o21ai_1
X_15601_ _06479_ _06481_ _09199_ _09581_ VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__o2bb2ai_2
X_12813_ _03636_ _03641_ _03640_ VGND VGND VPWR VPWR _03742_ sky130_fd_sc_hd__o21ai_1
X_13793_ _04585_ _04683_ net211 _04563_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a31oi_4
XFILLER_28_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15532_ net627 net532 net528 net631 VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__a22o_1
X_18320_ _09164_ _09160_ _09133_ _09165_ VGND VGND VPWR VPWR _09169_ sky130_fd_sc_hd__o211a_1
X_12744_ net645 net504 _03672_ _03673_ VGND VGND VPWR VPWR _03674_ sky130_fd_sc_hd__a22o_1
X_18251_ _09019_ _09097_ VGND VGND VPWR VPWR _09098_ sky130_fd_sc_hd__nand2_1
X_12675_ _03491_ _03370_ _03494_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__o21ai_1
X_17202_ net1093 _07924_ net503 _07926_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__a31o_1
X_15463_ _09384_ _09515_ _06350_ _06352_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__o22a_1
X_11626_ _02564_ _02560_ _02563_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__a21oi_2
X_18182_ _09026_ _09027_ VGND VGND VPWR VPWR _09029_ sky130_fd_sc_hd__nand2_1
X_15394_ net716 _06281_ _06282_ net657 _06277_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_41_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _05312_ _05313_ _05315_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__and3_1
XFILLER_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _08000_ _07895_ _07999_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__nand3b_1
X_11557_ net658 net535 VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__and2_1
XFILLER_7_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14345_ _05107_ _05247_ _05248_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__nand3_2
X_10508_ term_high\[56\] _01660_ net796 VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__a21oi_1
Xwire584 a_l\[9\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__buf_12
XFILLER_116_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap306 _08829_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__buf_1
X_17064_ _07930_ _07822_ VGND VGND VPWR VPWR _07933_ sky130_fd_sc_hd__nand2_1
XFILLER_7_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap317 _04937_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_2
XFILLER_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11488_ _02423_ _02424_ net269 VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__nand3_1
X_16015_ _06874_ _06875_ _06883_ _06884_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__o2bb2ai_2
Xmax_cap328 _01970_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__buf_4
Xmax_cap339 _08380_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_1
X_14276_ net315 _05141_ _05178_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__o21a_1
X_10439_ _01595_ _01599_ net443 _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__a31o_1
X_13227_ net796 _04142_ _04143_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__nor3_1
X_13158_ _04079_ _04058_ _04078_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__nor3_1
X_12109_ net698 net692 net483 net481 VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__nand4_2
X_17966_ net797 _08817_ _08818_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__nor3_1
XFILLER_88_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13089_ _04012_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__nand2_1
X_16917_ _07668_ _07784_ net1069 net503 _07783_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__o2111ai_2
XFILLER_78_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19705_ _00903_ _00905_ _00906_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__a21oi_2
XFILLER_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17897_ a_l\[14\] a_l\[15\] net480 net477 VGND VGND VPWR VPWR _08756_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_144_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16848_ _07713_ _07714_ _07589_ VGND VGND VPWR VPWR _07719_ sky130_fd_sc_hd__a21oi_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19636_ _00833_ _00832_ _00731_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__nand3_4
X_16779_ _07644_ _07647_ _07639_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__nand3_1
X_19567_ net367 _00756_ _00760_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__o21ai_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18518_ _09380_ _09382_ _09365_ VGND VGND VPWR VPWR _09385_ sky130_fd_sc_hd__a21o_1
X_19498_ _00490_ _00528_ _00529_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__nand3_1
X_18449_ _09187_ _09189_ _09304_ _09306_ VGND VGND VPWR VPWR _09310_ sky130_fd_sc_hd__o211ai_1
XFILLER_61_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20411_ clknet_leaf_30_clk _00051_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20342_ net793 net6 VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__and2_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20273_ _01512_ _01517_ _01516_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__a21o_1
XFILLER_1_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10790_ _01786_ _01810_ net405 VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__o21a_1
XFILLER_25_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12460_ _09624_ _03388_ _03383_ _03387_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__o211a_1
XFILLER_40_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11411_ _02349_ _02347_ net401 VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__and3_4
X_12391_ _03321_ _03323_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__nand2_1
X_20609_ clknet_leaf_35_clk _00249_ VGND VGND VPWR VPWR p_ll_pipe\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11342_ _09460_ _09592_ _01857_ _02278_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_49_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14130_ _05000_ _05005_ _05030_ _05004_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__o211ai_1
XFILLER_126_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11273_ _02185_ _02186_ _02208_ _02210_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_111_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14061_ _04964_ _04965_ _04966_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__a21oi_1
XFILLER_4_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10224_ net497 VGND VGND VPWR VPWR _09624_ sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_95_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13012_ _03857_ _03863_ _03933_ _03934_ VGND VGND VPWR VPWR _03939_ sky130_fd_sc_hd__nand4_1
X_17820_ _08680_ _08675_ _08679_ VGND VGND VPWR VPWR _08681_ sky130_fd_sc_hd__and3_1
XFILLER_79_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17751_ _08612_ _08613_ VGND VGND VPWR VPWR _08614_ sky130_fd_sc_hd__and2b_1
X_14963_ _05819_ _05820_ _05859_ _05860_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__nand4_1
X_16702_ _07443_ _07567_ _07568_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__nand3_2
X_17682_ _08544_ _08543_ VGND VGND VPWR VPWR _08546_ sky130_fd_sc_hd__nand2_1
XFILLER_75_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13914_ _04819_ _04812_ _04701_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__o211ai_4
X_14894_ _05707_ net263 _05743_ _05705_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_126_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16633_ _07497_ _07499_ _07494_ VGND VGND VPWR VPWR _07505_ sky130_fd_sc_hd__a21o_1
X_19421_ _09242_ _09308_ _04555_ _06985_ _00599_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__o221ai_2
X_13845_ _04747_ _04749_ _04743_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__a21oi_4
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19352_ _00524_ _00525_ _00527_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__a21o_1
X_16564_ _07302_ _07305_ _07306_ _07181_ _07182_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__o2111a_1
X_10988_ _01895_ _01905_ _01929_ _01930_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__o211ai_4
X_18303_ _09062_ _09148_ VGND VGND VPWR VPWR _09150_ sky130_fd_sc_hd__nand2_1
X_13776_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__inv_2
X_16495_ _07247_ _07250_ _07240_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__o21ai_1
X_15515_ net631 net627 VGND VGND VPWR VPWR _06401_ sky130_fd_sc_hd__and2_4
X_12727_ _03652_ _03653_ _03634_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__a21o_1
X_19283_ net754 net575 VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__nand2_1
X_12658_ _03576_ _03578_ _03587_ VGND VGND VPWR VPWR _03589_ sky130_fd_sc_hd__a21o_1
X_18234_ _09058_ _09075_ _08980_ VGND VGND VPWR VPWR _09081_ sky130_fd_sc_hd__a21boi_1
X_15446_ _06336_ net155 net795 _06337_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__o211a_1
X_11609_ _02546_ _02547_ _02476_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__a21o_1
X_18165_ _09011_ _09012_ VGND VGND VPWR VPWR _09013_ sky130_fd_sc_hd__nand2_1
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17116_ _07761_ _07768_ _07980_ _07981_ VGND VGND VPWR VPWR _07985_ sky130_fd_sc_hd__o22ai_1
Xclkbuf_leaf_10_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_12589_ _03512_ _03421_ _03511_ _03516_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__a31oi_1
X_15377_ net719 net649 _06267_ _06268_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__a22o_1
Xhold417 p_hh_pipe\[12\] VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold406 p_hh_pipe\[28\] VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18096_ _08887_ _08831_ _08885_ VGND VGND VPWR VPWR _08945_ sky130_fd_sc_hd__a21oi_2
Xwire370 _09505_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_1
X_14328_ _05223_ _05224_ _05226_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__a21oi_1
Xhold428 mid_sum\[24\] VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap147 _02811_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17047_ _07646_ _07814_ _07911_ _07913_ VGND VGND VPWR VPWR _07916_ sky130_fd_sc_hd__o211ai_4
Xhold439 p_ll\[11\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap158 _01540_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_1
X_14259_ net788 net783 net639 net636 VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__nand4_4
XFILLER_98_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _09883_ _09882_ _09887_ VGND VGND VPWR VPWR _09889_ sky130_fd_sc_hd__o21ai_4
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17949_ _08776_ _08804_ VGND VGND VPWR VPWR _08806_ sky130_fd_sc_hd__nand2_1
XFILLER_78_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19619_ _00809_ _00813_ _00782_ _00814_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__o211a_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20325_ net793 net22 VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__and2_1
XFILLER_134_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap681 net682 VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__buf_12
Xmax_cap670 net861 VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__buf_8
X_20256_ _01447_ _01488_ _01495_ _01454_ _01487_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__a221o_1
XFILLER_143_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20187_ net1013 net728 net557 net1096 _01376_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__a41o_1
X_11960_ net633 net546 VGND VGND VPWR VPWR _02896_ sky130_fd_sc_hd__nand2_1
X_10911_ net710 net704 VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nand2_8
XFILLER_45_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11891_ net698 net483 net481 net706 VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__a22o_1
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10842_ net795 net1182 VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__and2_1
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13630_ _04511_ _04512_ _04535_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__o21ai_2
X_10773_ _01792_ _01793_ _01797_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__nor3_1
X_13561_ _04320_ _04368_ _04369_ _04372_ _04266_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__a32oi_2
XFILLER_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16280_ _07151_ _07150_ _07090_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__nand3_4
X_12512_ net354 _03440_ _03443_ VGND VGND VPWR VPWR _03444_ sky130_fd_sc_hd__a21oi_1
XFILLER_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15300_ _06119_ _06123_ _06192_ _06108_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_57_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13492_ net768 net683 VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__nand2_1
XFILLER_12_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15231_ _06122_ _06123_ _06090_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__nand3_4
X_12443_ _03372_ _03374_ _03375_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_97_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12374_ _03187_ _03188_ _03185_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a21o_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15162_ _05989_ _06057_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__nand2_1
XFILLER_126_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11325_ _02265_ _02264_ _02263_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__nand3b_1
X_19970_ _01143_ _01149_ _01190_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__nand3_2
X_15093_ _05920_ _05955_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__nand2_1
X_14113_ _09264_ _09439_ _05013_ _05014_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__o211ai_4
XFILLER_140_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11256_ _02192_ _02194_ _02189_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__a21o_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18921_ net792 net553 VGND VGND VPWR VPWR _09813_ sky130_fd_sc_hd__nand2_1
X_14044_ _04945_ _04947_ _04869_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__a21bo_1
X_11187_ _02040_ _02041_ _02126_ _02128_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_128_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_66_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10207_ net998 VGND VGND VPWR VPWR _09439_ sky130_fd_sc_hd__clkinv_8
X_18852_ net621 net889 net1043 net1099 VGND VGND VPWR VPWR _09744_ sky130_fd_sc_hd__nand4_2
X_15995_ net1070 _06867_ net583 net541 _06865_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__o2111ai_4
XFILLER_94_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17803_ _08628_ _08662_ _08663_ VGND VGND VPWR VPWR _08665_ sky130_fd_sc_hd__nand3b_1
XFILLER_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18783_ _09670_ _09651_ VGND VGND VPWR VPWR _09674_ sky130_fd_sc_hd__nand2_1
X_17734_ _02589_ _07234_ _08486_ _08511_ _08517_ VGND VGND VPWR VPWR _08597_ sky130_fd_sc_hd__o2111ai_4
X_14946_ _05833_ _05834_ _05840_ _05841_ VGND VGND VPWR VPWR _05845_ sky130_fd_sc_hd__o2bb2ai_1
Xclkbuf_leaf_59_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_141_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17665_ _08523_ _08525_ _08478_ VGND VGND VPWR VPWR _08529_ sky130_fd_sc_hd__o21ai_1
X_14877_ _05771_ _05772_ net163 _05655_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__o211ai_2
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16616_ _07483_ _07484_ _07485_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_106_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ _08269_ _08270_ _08366_ _08367_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__and4_1
X_13828_ net762 net676 VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__nand2_1
X_19404_ _00583_ _00585_ _00580_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__a21oi_2
X_16547_ _07344_ _07346_ _07415_ _07416_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__a22o_1
X_13759_ _04665_ net432 net714 net963 _04554_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_18_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19335_ _05044_ _06605_ net618 net718 _00510_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__o2111ai_4
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_75_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19266_ b_l\[3\] net552 VGND VGND VPWR VPWR _10167_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16478_ _07256_ _07279_ _07257_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__a21boi_1
X_18217_ net791 net585 VGND VGND VPWR VPWR _09064_ sky130_fd_sc_hd__nand2_1
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19197_ _04555_ _06761_ _10086_ VGND VGND VPWR VPWR _10093_ sky130_fd_sc_hd__o21ai_2
X_15429_ _06275_ _06317_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__nand2_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18148_ _08980_ _08982_ _08992_ _08993_ VGND VGND VPWR VPWR _08996_ sky130_fd_sc_hd__o2bb2ai_1
X_18079_ _08924_ _08914_ _08923_ VGND VGND VPWR VPWR _08928_ sky130_fd_sc_hd__nand3_2
XFILLER_116_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20110_ _01270_ net143 _01179_ _01181_ _01269_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__o2111ai_4
XPHY_EDGE_ROW_84_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20041_ _01270_ net143 VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__nor2_1
XFILLER_112_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer311 b_h\[2\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer322 _09030_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__buf_1
XFILLER_10_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer300 net1095 VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer333 _04487_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer355 net1149 VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__buf_1
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11110_ _02053_ _01984_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__nand2_1
XFILLER_108_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20308_ _01552_ _01548_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__nand2_1
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12090_ net323 _02891_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_92_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11041_ _01984_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__nor2_2
X_20239_ _01480_ _01481_ net250 VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__a21oi_1
X_14800_ _05569_ _05572_ _05575_ _05692_ _05693_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__o2111ai_1
X_15780_ _06577_ _06658_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__nand2_2
X_12992_ _03913_ _03915_ _03900_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__o21ai_1
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11943_ _02708_ net438 _02873_ net358 VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__o211ai_1
X_14731_ _05630_ _05621_ _05601_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__o211ai_4
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11874_ _02693_ _02807_ _02808_ _02809_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__o31ai_2
X_17450_ net448 _08314_ _08302_ _08315_ VGND VGND VPWR VPWR _08316_ sky130_fd_sc_hd__o211a_2
XFILLER_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14662_ _04988_ _05285_ _05452_ _05560_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__o211ai_1
X_16401_ _07270_ _07272_ _07258_ VGND VGND VPWR VPWR _07275_ sky130_fd_sc_hd__a21oi_1
X_17381_ _08095_ _08099_ _08123_ _08126_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__o211ai_4
X_10825_ _01832_ _01839_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__and2_1
XFILLER_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13613_ net1058 net785 net666 net660 VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__nand4_4
X_16332_ _07199_ _07202_ net420 VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__a21o_1
XFILLER_60_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_861 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14593_ _05490_ _05491_ _05493_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__nand3_2
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19120_ _09910_ net1148 net592 net458 _06984_ VGND VGND VPWR VPWR _10010_ sky130_fd_sc_hd__a32o_1
X_10756_ _01756_ _01758_ _01783_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__a21boi_1
X_13544_ _04321_ _04324_ net352 _04451_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a22oi_1
X_16263_ _07000_ _07137_ _07136_ _07133_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_101_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13475_ _04384_ _04385_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__and2_1
X_10687_ _01723_ _01724_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__and2b_1
XFILLER_13_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19051_ net808 net562 VGND VGND VPWR VPWR _09942_ sky130_fd_sc_hd__nand2_1
X_16194_ _02338_ _06480_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__nor2_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12426_ _03346_ _03347_ _03354_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__a21o_1
X_18002_ _08834_ _08847_ _08852_ VGND VGND VPWR VPWR _08853_ sky130_fd_sc_hd__o21ai_2
X_15214_ _06009_ _06107_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__nand2_1
X_15145_ _06037_ _06040_ _06005_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_134_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12357_ _03273_ _03275_ _03288_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__nand3_2
X_11308_ _02246_ _02247_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__nand2_2
X_12288_ _03038_ _03064_ _03065_ _03069_ _03072_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__a32oi_4
XFILLER_107_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19953_ _01166_ _01168_ _01171_ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__a21o_1
X_15076_ _05967_ _05969_ _05902_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__o21ai_1
X_11239_ _02161_ _02162_ _02178_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o21ai_1
X_18904_ _09669_ _09795_ VGND VGND VPWR VPWR _09796_ sky130_fd_sc_hd__nand2_1
X_19884_ net894 net1102 net548 net820 VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__a22oi_2
X_14027_ _04931_ _04920_ _04930_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__nand3_2
X_18835_ _09725_ _09727_ _09582_ VGND VGND VPWR VPWR _09728_ sky130_fd_sc_hd__a21oi_2
XFILLER_83_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15978_ _06784_ net283 _06787_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__a21boi_2
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18766_ _09155_ _09297_ VGND VGND VPWR VPWR _09655_ sky130_fd_sc_hd__nor2_1
X_17717_ _08575_ _08576_ _08562_ VGND VGND VPWR VPWR _08580_ sky130_fd_sc_hd__a21oi_4
X_18697_ _09444_ _09578_ _09579_ VGND VGND VPWR VPWR _09580_ sky130_fd_sc_hd__nand3_2
X_14929_ net739 net733 net663 net655 _05826_ VGND VGND VPWR VPWR _05828_ sky130_fd_sc_hd__a41o_1
XFILLER_91_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17648_ _08381_ _08505_ _08506_ VGND VGND VPWR VPWR _08512_ sky130_fd_sc_hd__nand3_4
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17579_ _08438_ _08440_ _08429_ _08431_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__o211ai_1
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20590_ clknet_leaf_12_clk _00230_ VGND VGND VPWR VPWR p_hh_pipe\[20\] sky130_fd_sc_hd__dfxtp_1
X_19318_ _10010_ _10027_ _10026_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__a21boi_4
X_19249_ _09868_ _09988_ _09990_ _09737_ VGND VGND VPWR VPWR _10150_ sky130_fd_sc_hd__a31oi_4
XFILLER_129_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_132_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20024_ _01251_ _01252_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__nand2_1
XFILLER_132_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer51 _06401_ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__buf_4
Xrebuffer62 b_h\[9\] VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer40 a_h\[11\] VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer73 a_h\[12\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer84 b_l\[2\] VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer95 b_l\[4\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11590_ _02523_ _02525_ net692 net501 VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__nand4_4
X_20788_ clknet_leaf_7_clk _00428_ VGND VGND VPWR VPWR a_l\[10\] sky130_fd_sc_hd__dfxtp_4
X_10610_ net794 net1228 VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_12_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ net793 net1214 VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__and2_1
XFILLER_128_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer141 net936 VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd1_1
X_13260_ _04171_ _04172_ _04173_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__a21o_1
Xrebuffer130 _09889_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__buf_2
X_10472_ _01632_ net140 net793 _01633_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__o211a_1
Xrebuffer152 _02804_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlymetal6s4s_1
XFILLER_108_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12211_ _03138_ _03139_ _03141_ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__a21o_1
Xrebuffer174 net611 VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer163 a_l\[13\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer185 _02334_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer196 b_h\[7\] VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd1_1
X_13191_ _04112_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__inv_2
XFILLER_123_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ _03068_ net268 _03072_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__a21o_1
X_16950_ net558 net523 net516 net566 VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__a22o_1
X_12073_ net644 net526 VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__nand2_2
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15901_ _09199_ _09602_ _06774_ _06775_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__o211ai_2
X_11024_ _01957_ _01966_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__nand2_2
XFILLER_89_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16881_ net586 net498 VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__nand2_1
XFILLER_89_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15832_ _06709_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__nand2_2
XFILLER_66_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18620_ _09488_ _09490_ _09477_ VGND VGND VPWR VPWR _09496_ sky130_fd_sc_hd__nand3_4
XFILLER_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15763_ _06560_ _06563_ _06638_ _06639_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__o211ai_2
X_18551_ _09416_ _09418_ VGND VGND VPWR VPWR _09421_ sky130_fd_sc_hd__and2b_1
XFILLER_58_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12975_ net645 net885 VGND VGND VPWR VPWR _03902_ sky130_fd_sc_hd__nand2_1
X_17502_ _08366_ _08367_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__nand2_1
X_11926_ net665 net511 VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__nand2_4
X_18482_ net801 net610 net458 _09269_ _09274_ VGND VGND VPWR VPWR _09345_ sky130_fd_sc_hd__a32o_1
X_14714_ net736 net670 net668 net740 VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__a22o_1
XFILLER_17_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _06573_ _06574_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__nor2_1
X_17433_ _08221_ _08227_ _08295_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__o21ai_2
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11857_ _02788_ _02789_ _02791_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__nand3_1
X_14645_ _05544_ _05545_ _05541_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__a21o_1
X_10808_ _01828_ _01827_ net796 VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__a21oi_1
X_11788_ net652 net1023 VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__nand2_1
X_17364_ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__inv_2
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14576_ net730 net685 VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16315_ _02338_ _06480_ _07066_ _07067_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_136_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17295_ _08161_ _08162_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__nor2_1
X_10739_ p_hl\[16\] p_lh\[16\] p_hl\[17\] p_lh\[17\] VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__a22o_1
X_13527_ _04434_ _04436_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__nand2_1
X_19103_ _09988_ _09990_ _09868_ VGND VGND VPWR VPWR _09994_ sky130_fd_sc_hd__a21oi_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16246_ _07108_ _07119_ _07109_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__nand3_2
X_19034_ _09808_ _09826_ _09823_ _09820_ VGND VGND VPWR VPWR _09925_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_146_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13458_ _04367_ _04333_ VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__nand2_1
Xoutput105 net105 VGND VGND VPWR VPWR p[45] sky130_fd_sc_hd__buf_2
Xoutput116 net116 VGND VGND VPWR VPWR p[55] sky130_fd_sc_hd__buf_2
X_16177_ _07051_ _07052_ _06949_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__a21oi_4
XFILLER_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12409_ _03299_ _03337_ _03339_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__nand3_1
X_13389_ _04297_ _04298_ _04269_ VGND VGND VPWR VPWR _04301_ sky130_fd_sc_hd__a21oi_1
Xoutput127 net127 VGND VGND VPWR VPWR p[7] sky130_fd_sc_hd__buf_2
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15128_ _06023_ net657 net730 _06021_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__nand4_1
XFILLER_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19936_ _01158_ VGND VGND VPWR VPWR _01159_ sky130_fd_sc_hd__inv_2
X_15059_ _05936_ _05953_ _05954_ _05921_ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_56_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19867_ _01081_ _01082_ _01083_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_147_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18818_ _09709_ _09634_ VGND VGND VPWR VPWR _09711_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19798_ net591 net718 _01007_ _01008_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__a22oi_4
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18749_ net301 _09508_ _09495_ _09489_ VGND VGND VPWR VPWR _09637_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_36_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20711_ clknet_leaf_40_clk _00351_ VGND VGND VPWR VPWR p_lh\[13\] sky130_fd_sc_hd__dfxtp_1
X_20642_ clknet_leaf_18_clk _00282_ VGND VGND VPWR VPWR p_hh\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20573_ clknet_leaf_28_clk _00213_ VGND VGND VPWR VPWR p_hh_pipe\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20007_ _01232_ _01215_ _01233_ VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__and3_1
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_87_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _03686_ _03688_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__nand2_2
XFILLER_70_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11711_ net679 net508 VGND VGND VPWR VPWR _02649_ sky130_fd_sc_hd__nand2_1
X_12691_ _03618_ _03619_ net682 net474 VGND VGND VPWR VPWR _03621_ sky130_fd_sc_hd__nand4_2
X_11642_ _01888_ _02338_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__nor2_1
XFILLER_70_775 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14430_ net723 net695 VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__nand2_1
X_14361_ _05107_ _05247_ _05248_ _05089_ _05252_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__a32oi_4
X_16100_ _06875_ _06887_ _06874_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__a21boi_1
X_11573_ _02505_ _02507_ _02494_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__nand3_2
X_13312_ _04195_ _04222_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__nand2_1
Xwire711 a_h\[1\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__buf_12
XPHY_EDGE_ROW_30_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 a[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
X_10524_ net1355 _01669_ net1323 VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__a21oi_1
Xinput29 a[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17080_ _07749_ _07752_ _07755_ VGND VGND VPWR VPWR _07949_ sky130_fd_sc_hd__o21ai_2
XFILLER_7_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14292_ b_l\[14\] net709 _05192_ _05193_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__a22oi_2
Xwire744 net835 VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__buf_12
X_10455_ net793 _01618_ _01619_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__and3_1
X_16031_ _06903_ _06896_ _06904_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__nand3_4
XFILLER_109_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13243_ a_h\[0\] net766 net710 net923 VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__a22oi_1
XFILLER_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13174_ net320 _04074_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__or2_1
X_10386_ _01554_ _01559_ net796 VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__a21oi_1
X_12125_ net461 _03056_ _03048_ _03057_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__o211a_1
XFILLER_123_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17982_ _08831_ _08832_ VGND VGND VPWR VPWR _08833_ sky130_fd_sc_hd__nor2_1
XFILLER_78_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12056_ _02986_ _02988_ _02989_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__a21oi_2
X_16933_ _07793_ _07795_ _07799_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__o21ai_1
X_19721_ _09275_ _09308_ _00916_ _09297_ _00919_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__o221ai_2
X_11007_ net707 net517 _01947_ _01949_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__a22o_1
X_16864_ _07624_ _07625_ _07696_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__o21ai_1
X_19652_ _00702_ _00845_ _00847_ _00850_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__nand4_2
X_15815_ net587 net543 VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__nand2_1
X_18603_ _09369_ _09372_ _09375_ VGND VGND VPWR VPWR _09477_ sky130_fd_sc_hd__o21ai_2
X_16795_ _07512_ _07516_ _07514_ VGND VGND VPWR VPWR _07666_ sky130_fd_sc_hd__a21oi_2
X_19583_ net1074 _00770_ _00771_ _00775_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__nand4_2
X_15746_ _06586_ _06618_ _06619_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__nand3_1
XFILLER_73_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18534_ _09396_ _09387_ _09326_ _09398_ VGND VGND VPWR VPWR _09402_ sky130_fd_sc_hd__o211ai_4
X_12958_ net944 net474 _03881_ _03882_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a22o_1
X_11909_ _02832_ _02839_ _02840_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__nand3_1
X_15677_ _06552_ _06549_ _06510_ _06555_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__o211ai_1
X_18465_ _09265_ _09289_ _09266_ VGND VGND VPWR VPWR _09326_ sky130_fd_sc_hd__a21boi_4
X_12889_ net944 net478 _03812_ _03813_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__a22o_1
X_17416_ net795 _08281_ _08282_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__and3_1
X_18396_ net1123 net1146 net599 net593 VGND VGND VPWR VPWR _09251_ sky130_fd_sc_hd__nand4_4
X_14628_ _05384_ _05525_ _05524_ _05523_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__o211ai_1
X_17347_ _08052_ _08210_ _08206_ _08208_ VGND VGND VPWR VPWR _08214_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_44_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14559_ _05433_ _05434_ _05456_ _05458_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__nand4_2
XFILLER_147_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17278_ net160 _08003_ _08143_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__o21ai_2
X_16229_ _07099_ _07102_ _09297_ _09581_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__o2bb2ai_1
X_19017_ net753 net589 VGND VGND VPWR VPWR _09908_ sky130_fd_sc_hd__nand2_1
XFILLER_127_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19919_ _01130_ _01131_ net332 _01124_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__o211ai_2
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20625_ clknet_leaf_47_clk _00265_ VGND VGND VPWR VPWR p_ll_pipe\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20556_ clknet_leaf_18_clk _00196_ VGND VGND VPWR VPWR mid_sum\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10240_ net794 net64 VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__and2_1
X_20487_ clknet_leaf_45_clk _00127_ VGND VGND VPWR VPWR term_mid\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13930_ net714 net724 net709 net728 VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__a22oi_2
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15600_ _06479_ _06481_ _09199_ _09581_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__o2bb2a_1
X_13861_ _04767_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__inv_2
X_16580_ _07348_ _07416_ _07414_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__a21o_1
XFILLER_90_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12812_ _03739_ _03740_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__nor2_1
X_13792_ net796 _04698_ _04699_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__nor3b_1
X_15531_ net627 net532 net528 net631 VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__a22oi_1
X_12743_ net638 net634 b_h\[6\] net994 VGND VGND VPWR VPWR _03673_ sky130_fd_sc_hd__nand4_2
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18250_ net187 _09094_ _09095_ VGND VGND VPWR VPWR _09097_ sky130_fd_sc_hd__a21o_1
XFILLER_63_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15462_ _06350_ _06351_ net716 net643 VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__and4b_1
X_12674_ _03121_ _03603_ _03604_ _03117_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__nand4_4
X_17201_ _07921_ _07926_ _07924_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__o21ai_2
X_14413_ _05312_ _05313_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__a21oi_2
X_11625_ _02440_ _02561_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__nor2_1
X_18181_ net623 net626 net759 net754 VGND VGND VPWR VPWR _09028_ sky130_fd_sc_hd__nand4_2
X_15393_ _06283_ _06285_ _06277_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_41_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17132_ _07998_ _08000_ _07895_ VGND VGND VPWR VPWR _08001_ sky130_fd_sc_hd__o21bai_1
Xwire541 net903 VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__buf_12
X_11556_ _02364_ _02357_ _02360_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__a21oi_2
X_14344_ _05245_ _05242_ _05116_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__a21o_1
X_10507_ net796 _01659_ _01660_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__nor3_1
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap307 _07387_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__buf_6
X_17063_ _07924_ _07927_ _07922_ VGND VGND VPWR VPWR _07932_ sky130_fd_sc_hd__a21o_1
X_14275_ _05144_ net931 VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__nand2_1
X_11487_ _02424_ _02354_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__nand2_1
X_16014_ _06885_ _06886_ _06874_ _06875_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__o211ai_2
X_13226_ _04141_ _04133_ net710 net713 VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__and4_1
Xmax_cap329 _01418_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
X_10438_ term_mid\[41\] term_high\[41\] _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__o21a_1
XFILLER_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13157_ _04078_ _04079_ _04058_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__o21ai_1
X_10369_ term_low\[31\] term_mid\[31\] term_low\[30\] term_mid\[30\] VGND VGND VPWR
+ VPWR _01428_ sky130_fd_sc_hd__o211a_1
XFILLER_112_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12108_ net692 net481 VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__nand2_1
X_17965_ _08815_ _08816_ net459 _06402_ VGND VGND VPWR VPWR _08818_ sky130_fd_sc_hd__a211oi_1
XFILLER_69_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13088_ _03969_ _03968_ _04009_ _04008_ _04010_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__o2111ai_2
X_12039_ _09460_ _09613_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__nor2_1
X_16916_ net572 net570 net513 net506 VGND VGND VPWR VPWR _07786_ sky130_fd_sc_hd__nand4_2
X_19704_ _00903_ _00905_ _00906_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__and3_1
X_17896_ a_l\[15\] net480 net477 net555 VGND VGND VPWR VPWR _08755_ sky130_fd_sc_hd__a22o_1
XFILLER_93_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_144_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16847_ _07589_ _07713_ _07714_ VGND VGND VPWR VPWR _07718_ sky130_fd_sc_hd__nand3_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19635_ _00778_ _00831_ _00830_ _00732_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__o211ai_2
X_16778_ _07644_ _07647_ _07639_ VGND VGND VPWR VPWR _07649_ sky130_fd_sc_hd__a21o_1
X_19566_ _00750_ _00751_ _00739_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__nand3_4
XFILLER_19_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15729_ _06604_ _06607_ _06599_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__a21oi_1
X_18517_ _09365_ _09380_ _09382_ VGND VGND VPWR VPWR _09383_ sky130_fd_sc_hd__nand3_2
XFILLER_34_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19497_ _00635_ _00683_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__nand2_1
X_18448_ _09304_ _09190_ VGND VGND VPWR VPWR _09309_ sky130_fd_sc_hd__nand2_1
X_18379_ _09151_ _09154_ _09149_ VGND VGND VPWR VPWR _09233_ sky130_fd_sc_hd__a21oi_4
X_20410_ clknet_leaf_30_clk _00050_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfxtp_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20341_ net793 net5 VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__and2_1
XFILLER_115_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20272_ _01514_ _01515_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__nand2_1
XFILLER_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11410_ _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__inv_2
X_20608_ clknet_leaf_32_clk _00248_ VGND VGND VPWR VPWR p_ll_pipe\[6\] sky130_fd_sc_hd__dfxtp_1
X_12390_ _03317_ net460 _03308_ _03316_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__o211ai_2
XFILLER_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11341_ _02277_ _02279_ _02274_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a21o_1
XFILLER_20_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_104_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20539_ clknet_leaf_42_clk _00179_ VGND VGND VPWR VPWR mid_sum\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_4_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11272_ _02185_ _02186_ _02209_ _02211_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__nand4_1
X_14060_ _04964_ _04965_ _09690_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_111_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10223_ net504 VGND VGND VPWR VPWR _09613_ sky130_fd_sc_hd__inv_16
X_13011_ net175 _03935_ _03936_ _03937_ VGND VGND VPWR VPWR _03938_ sky130_fd_sc_hd__nand4_2
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17750_ _08611_ _08610_ _08609_ VGND VGND VPWR VPWR _08613_ sky130_fd_sc_hd__nand3_1
XFILLER_87_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14962_ _05819_ _05820_ _05859_ _05860_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__a22o_1
X_16701_ _07442_ _07570_ _07571_ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_113_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17681_ _08372_ _08452_ _08455_ _08543_ VGND VGND VPWR VPWR _08545_ sky130_fd_sc_hd__a31o_1
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13913_ _04814_ _04673_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__nand2_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14893_ _05707_ _05743_ net263 _05705_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_126_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16632_ _09242_ _09613_ _07353_ _07498_ _07497_ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__o221ai_4
XFILLER_90_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19420_ _00598_ _00600_ _00595_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__o21ai_2
X_13844_ _02502_ _04134_ net778 net660 _04747_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__o2111ai_4
XFILLER_90_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19351_ _00524_ _00525_ _00526_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__nand3_1
X_16563_ _07051_ _07177_ _07178_ _07304_ VGND VGND VPWR VPWR _07436_ sky130_fd_sc_hd__a211oi_2
X_10987_ _01906_ _01931_ _01932_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__nand3_1
X_18302_ net782 net585 net582 net791 VGND VGND VPWR VPWR _09149_ sky130_fd_sc_hd__a22oi_2
XFILLER_50_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13775_ _04682_ _04655_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__nand2_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16494_ _07365_ _07366_ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__nand2_1
X_15514_ _09690_ net1105 net631 VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__and3_1
X_12726_ _03630_ _03632_ _03652_ _03653_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__o211ai_2
X_19282_ net878 net567 VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__nand2_4
X_12657_ _03576_ _03578_ _03587_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18233_ _08973_ _08974_ _08978_ _08994_ VGND VGND VPWR VPWR _09080_ sky130_fd_sc_hd__a31o_1
X_15445_ net155 _06308_ net162 VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_122_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11608_ _02479_ _02543_ _02544_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__nand3_4
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18164_ _08953_ _08934_ _09008_ _09009_ VGND VGND VPWR VPWR _09012_ sky130_fd_sc_hd__o211ai_4
X_15376_ _06221_ _06264_ net719 net649 _06268_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__o2111ai_4
XFILLER_117_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17115_ _07746_ _07761_ _07760_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__o21ai_2
X_12588_ _09504_ _03510_ _03421_ _03512_ VGND VGND VPWR VPWR _03519_ sky130_fd_sc_hd__o211ai_2
XFILLER_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14327_ _05225_ _05226_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__nand2_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold407 p_hh_pipe\[13\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_129_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire382 _06609_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_2
X_11539_ _02383_ _02384_ net327 _02390_ _02416_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__a32oi_2
X_18095_ _08887_ _08831_ _08885_ VGND VGND VPWR VPWR _08944_ sky130_fd_sc_hd__a21o_1
Xhold418 mid_sum\[9\] VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 p_hh_pipe\[10\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17046_ _07646_ _07814_ _07911_ _07913_ VGND VGND VPWR VPWR _07915_ sky130_fd_sc_hd__o211a_1
X_14258_ net783 net636 VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__nand2_1
XFILLER_131_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13209_ _04127_ _04121_ VGND VGND VPWR VPWR _04130_ sky130_fd_sc_hd__nand2_1
X_14189_ _05084_ _05086_ _05091_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_51_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _09885_ _09886_ _09887_ VGND VGND VPWR VPWR _09888_ sky130_fd_sc_hd__a21o_1
XFILLER_100_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17948_ _08770_ _08791_ VGND VGND VPWR VPWR _08805_ sky130_fd_sc_hd__or2_1
XFILLER_39_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17879_ _08736_ _08737_ _08738_ VGND VGND VPWR VPWR _08739_ sky130_fd_sc_hd__o21ai_1
Xclone272 net1071 VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__clkbuf_16
Xclone261 net1087 VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__clkbuf_16
X_19618_ _00783_ _00815_ _00816_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__nand3_2
XFILLER_19_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19549_ b_l\[8\] net567 VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__nand2_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20324_ net793 net21 VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__and2_1
XFILLER_135_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap671 net672 VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__buf_8
X_20255_ _01447_ _01488_ _01495_ _01454_ _01487_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__a221oi_1
Xmax_cap660 net1025 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__buf_8
XFILLER_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap682 net684 VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__buf_12
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20186_ _09297_ _09384_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__nor2_1
XFILLER_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10910_ net713 net1106 VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__nand2_1
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_450 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11890_ _02701_ _02715_ _02714_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__o21a_1
X_10841_ net795 net1322 VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_121_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10772_ net442 _01785_ _01789_ _01796_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__a31o_1
XFILLER_71_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13560_ _04371_ _04319_ _04370_ _04265_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__a31oi_1
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12511_ net1019 _03260_ b_h\[8\] _03262_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__a31o_1
X_13491_ net763 net694 VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__nand2_1
X_12442_ _03372_ _03374_ net793 VGND VGND VPWR VPWR _03375_ sky130_fd_sc_hd__o21ai_1
XFILLER_9_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15230_ _06090_ _06124_ _06125_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_97_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12373_ _03304_ _03305_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15161_ _06053_ _05988_ _06052_ VGND VGND VPWR VPWR _06058_ sky130_fd_sc_hd__nand3_2
X_11324_ _02189_ _02194_ _02191_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15092_ _05902_ _05968_ _05969_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__a21oi_2
X_14112_ _05014_ _05013_ _05011_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__a21o_1
X_11255_ _02104_ _02193_ _02189_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__o21ai_2
X_18920_ net1064 net557 VGND VGND VPWR VPWR _09812_ sky130_fd_sc_hd__nand2_1
X_14043_ _04945_ _04947_ _04869_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__a21o_1
XFILLER_140_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10206_ a_h\[5\] VGND VGND VPWR VPWR _09428_ sky130_fd_sc_hd__inv_12
X_11186_ _02126_ _02128_ _02043_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18851_ net621 net1043 net1099 net889 VGND VGND VPWR VPWR _09743_ sky130_fd_sc_hd__a22o_1
X_15994_ _06864_ _06868_ _06861_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__o21bai_1
X_17802_ _08662_ _08663_ _08628_ VGND VGND VPWR VPWR _08664_ sky130_fd_sc_hd__a21bo_1
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18782_ _09647_ _09648_ _09667_ _09669_ VGND VGND VPWR VPWR _09673_ sky130_fd_sc_hd__o211ai_1
X_17733_ _08482_ _08485_ _08595_ VGND VGND VPWR VPWR _08596_ sky130_fd_sc_hd__o21ai_2
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14945_ _05840_ _05841_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17664_ _08474_ _08476_ _08524_ _08526_ VGND VGND VPWR VPWR _08528_ sky130_fd_sc_hd__o211ai_1
X_14876_ _05771_ _05772_ net163 _05655_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__o211a_1
X_19403_ _05044_ _06605_ _00512_ _00525_ _00582_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__o2111ai_4
X_16615_ _07484_ _07485_ VGND VGND VPWR VPWR _07487_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_106_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17595_ _08270_ _08367_ _08365_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__a21oi_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13827_ net773 net1122 net670 net667 VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__nand4_4
X_16546_ _07348_ _07416_ VGND VGND VPWR VPWR _07419_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13758_ _04663_ _04664_ _04661_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__a21oi_1
XFILLER_16_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19334_ _05044_ _06605_ net618 net718 _00510_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__o2111a_1
X_12709_ net654 net648 net859 VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__nand3_2
X_19265_ net919 net556 VGND VGND VPWR VPWR _10166_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_139_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16477_ _07257_ _07349_ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__nand2_1
XFILLER_86_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18216_ net782 net593 VGND VGND VPWR VPWR _09063_ sky130_fd_sc_hd__nand2_1
X_13689_ net789 net785 net660 net656 VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_61_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19196_ _10089_ _10091_ _10086_ VGND VGND VPWR VPWR _10092_ sky130_fd_sc_hd__a21oi_4
X_15428_ _06274_ _06318_ _06271_ _06272_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__nand4_1
X_18147_ _08989_ _08991_ _08972_ _08981_ _08980_ VGND VGND VPWR VPWR _08995_ sky130_fd_sc_hd__o221ai_2
X_15359_ _06249_ _06250_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__o21bai_2
XFILLER_144_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18078_ _08924_ _08914_ VGND VGND VPWR VPWR _08927_ sky130_fd_sc_hd__nand2_2
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17029_ net978 _07808_ _07813_ _07824_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__a31oi_4
X_20040_ net203 _01264_ _01174_ _01167_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer312 net530 VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__buf_6
Xrebuffer301 net1095 VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_79_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer334 net770 VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20307_ _01546_ net152 _01551_ _01502_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__o22ai_1
XFILLER_146_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap490 b_h\[11\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_12
XFILLER_1_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11040_ _01982_ _01983_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__and2_1
XFILLER_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20238_ _09297_ _09384_ _01429_ _01431_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__o31ai_2
XFILLER_130_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20169_ net735 net551 _09308_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__a21o_1
X_12991_ _03896_ _03898_ _03913_ _03915_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_123_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11942_ _02708_ net438 _02873_ _02872_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__o211a_1
XFILLER_55_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14730_ _05622_ _05625_ _05608_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__a21o_1
XFILLER_18_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11873_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__inv_2
XFILLER_55_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14661_ _05561_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__inv_2
X_16400_ _07258_ _07270_ _07272_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__nand3_1
X_17380_ _08124_ _08245_ _08246_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__nand3_1
X_10824_ p_hl\[30\] net1366 VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__xnor2_1
X_13612_ _04416_ _04519_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__nand2_1
X_14592_ _05488_ _05492_ _05489_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__nand3_2
XFILLER_32_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16331_ net629 a_l\[0\] _02588_ _07203_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__a31o_1
X_13543_ _04438_ net352 _04451_ VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__nand3_2
XFILLER_13_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10755_ _01754_ _01762_ _01767_ _01774_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__and4b_1
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16262_ _06996_ _06997_ _06995_ VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_101_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13474_ _04314_ _04317_ _04383_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__a21o_1
X_10686_ p_hl\[10\] p_lh\[10\] VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__nand2_2
X_19050_ net1146 net568 net1084 net775 VGND VGND VPWR VPWR _09941_ sky130_fd_sc_hd__a22o_1
XFILLER_145_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16193_ net620 net496 net491 net841 VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__a22o_1
X_12425_ _03346_ _03347_ _03354_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__nand3_1
X_18001_ _08834_ _08847_ _08850_ _08826_ VGND VGND VPWR VPWR _08852_ sky130_fd_sc_hd__a22oi_1
X_15213_ net726 net722 a_h\[10\] net657 VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__nand4_1
X_12356_ _03287_ _03288_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__nand2_1
X_15144_ _06040_ _06005_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_134_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11307_ _02246_ _02247_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__and2_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ net698 net692 net463 _03045_ VGND VGND VPWR VPWR _03221_ sky130_fd_sc_hd__a31oi_4
X_19952_ _01059_ _01166_ _01168_ _01169_ VGND VGND VPWR VPWR _01177_ sky130_fd_sc_hd__nand4_2
XFILLER_4_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15075_ _05900_ _05901_ _05968_ _05970_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__nand4_1
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11238_ _02176_ _02177_ net362 VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__nand3_1
X_18903_ _09651_ _09667_ VGND VGND VPWR VPWR _09795_ sky130_fd_sc_hd__nand2_1
X_19883_ net820 net894 net1102 net548 VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__and4_2
X_14026_ _04921_ _04928_ _04929_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__nand3_2
X_11169_ _09177_ _09613_ _02106_ _02108_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__o211ai_1
XFILLER_68_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18834_ _09720_ _09722_ _09724_ VGND VGND VPWR VPWR _09727_ sky130_fd_sc_hd__nand3_1
XFILLER_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15977_ _06787_ _06817_ VGND VGND VPWR VPWR _06854_ sky130_fd_sc_hd__nand2_1
X_18765_ _09480_ _09653_ VGND VGND VPWR VPWR _09654_ sky130_fd_sc_hd__nand2_1
X_17716_ _08561_ _08575_ _08576_ VGND VGND VPWR VPWR _08579_ sky130_fd_sc_hd__nand3_1
X_18696_ _09575_ net275 VGND VGND VPWR VPWR _09579_ sky130_fd_sc_hd__nand2_1
X_14928_ _05824_ _05825_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17647_ _08509_ net339 _08508_ VGND VGND VPWR VPWR _08511_ sky130_fd_sc_hd__nand3_4
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14859_ _05754_ _05755_ _05757_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__a21o_1
XFILLER_24_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17578_ _08439_ _08441_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__nand2_1
XFILLER_51_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19317_ _10010_ _10027_ _10025_ _10020_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__o2bb2ai_4
X_16529_ net307 _07389_ _07399_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__nand3_1
X_19248_ _10140_ _10141_ _10143_ VGND VGND VPWR VPWR _10149_ sky130_fd_sc_hd__nand3_1
X_19179_ net369 _09890_ _09893_ VGND VGND VPWR VPWR _10074_ sky130_fd_sc_hd__a21o_1
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_104_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20023_ _01248_ _01246_ _01201_ VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nand3_4
XFILLER_132_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer30 net824 VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_27_623 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer52 net848 VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer63 _02495_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer41 a_h\[11\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer74 net870 VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer96 b_l\[8\] VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer85 b_l\[2\] VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlymetal6s2s_1
X_20787_ clknet_leaf_19_clk _00427_ VGND VGND VPWR VPWR a_l\[9\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_12_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ net793 net1235 VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__and2_1
XFILLER_22_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10471_ _01626_ _01630_ _01631_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__o21ai_1
Xrebuffer131 a_l\[5\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer120 net915 VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_136_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer142 net936 VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__buf_1
X_12210_ _03138_ _03139_ _03141_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__nand3_2
Xrebuffer164 net960 VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer175 a_l\[0\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer197 b_h\[7\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd1_1
X_13190_ _04105_ _04110_ _04109_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__a21bo_1
XFILLER_135_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12141_ _03072_ net268 _03068_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__nand3b_2
X_12072_ net644 net524 VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__nand2_2
X_15900_ _06771_ _06774_ _06775_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__and3_1
X_11023_ _01961_ _01963_ _01959_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__a21o_1
XFILLER_103_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16880_ net594 net493 VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__nand2_1
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15831_ _06673_ _06708_ _06707_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__nand3_2
X_15762_ _06638_ _06639_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__nand2_1
X_18550_ _09412_ _09413_ _09415_ VGND VGND VPWR VPWR _09420_ sky130_fd_sc_hd__and3_1
X_12974_ _03897_ _03899_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__nand2_1
X_11925_ _02753_ _02719_ _02752_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__a21boi_2
X_17501_ _08362_ _08363_ _08364_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__nand3_2
X_18481_ _09328_ _09339_ _09341_ VGND VGND VPWR VPWR _09344_ sky130_fd_sc_hd__nand3_2
X_14713_ net740 net668 VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__nand2_1
XFILLER_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _06504_ _06571_ _06572_ net797 VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__a31o_1
X_17432_ _08292_ _08294_ _08221_ _08227_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11856_ _02790_ _02792_ VGND VGND VPWR VPWR _02793_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14644_ _05333_ _05467_ _05472_ _05494_ _05500_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__o2111ai_4
X_11787_ _02628_ _02722_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__nand2_1
X_10807_ p_hl\[26\] net1306 _01826_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a21bo_1
X_17363_ _08077_ _08074_ _08048_ _08229_ VGND VGND VPWR VPWR _08230_ sky130_fd_sc_hd__o211ai_4
XFILLER_9_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14575_ _05343_ _05348_ _05345_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_31_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16314_ _02338_ _06480_ _07066_ _07067_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__o22ai_2
XTAP_TAPCELL_ROW_136_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17294_ _08020_ _08030_ _08160_ net796 VGND VGND VPWR VPWR _08162_ sky130_fd_sc_hd__a31o_1
X_10738_ _01754_ _01759_ _01762_ VGND VGND VPWR VPWR _01768_ sky130_fd_sc_hd__nand3b_1
X_13526_ _04400_ _04432_ _04433_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__nand3_1
X_19102_ _09976_ _09977_ _09987_ VGND VGND VPWR VPWR _09993_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_136_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16245_ _07111_ _07118_ _07116_ VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__o21ai_2
X_13457_ _04331_ _04332_ _04365_ _04366_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__nand4_2
X_19033_ _09922_ _09923_ VGND VGND VPWR VPWR _09924_ sky130_fd_sc_hd__nand2_4
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ _03295_ _03298_ _03334_ _03335_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__nand4_1
X_10669_ p_hl\[7\] p_lh\[7\] VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__or2_1
Xoutput106 net106 VGND VGND VPWR VPWR p[46] sky130_fd_sc_hd__buf_2
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16176_ net154 _07047_ _06950_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__a21o_4
X_13388_ _04294_ _04295_ _04280_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__a21o_1
Xoutput117 net117 VGND VGND VPWR VPWR p[56] sky130_fd_sc_hd__buf_2
Xoutput128 net128 VGND VGND VPWR VPWR p[8] sky130_fd_sc_hd__buf_2
X_12339_ _03268_ _03269_ _03253_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__a21oi_1
X_15127_ _06021_ _06023_ _09308_ _09493_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19935_ _01156_ _01155_ VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__nand2_2
X_15058_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__inv_2
XFILLER_141_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14009_ net351 _04872_ _04910_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__o21ai_2
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19866_ _01081_ _01082_ net794 VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18817_ _09632_ _09633_ _09707_ _09708_ VGND VGND VPWR VPWR _09710_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_39_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19797_ _01008_ net718 net591 _01007_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_39_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18748_ _09473_ _09512_ _09514_ _09517_ VGND VGND VPWR VPWR _09636_ sky130_fd_sc_hd__o2bb2ai_1
X_20710_ clknet_leaf_40_clk _00350_ VGND VGND VPWR VPWR p_lh\[12\] sky130_fd_sc_hd__dfxtp_1
X_18679_ _09412_ _09553_ _09555_ VGND VGND VPWR VPWR _09561_ sky130_fd_sc_hd__nand3_1
XFILLER_51_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20641_ clknet_leaf_18_clk _00281_ VGND VGND VPWR VPWR p_hh\[7\] sky130_fd_sc_hd__dfxtp_1
X_20572_ clknet_leaf_26_clk _00212_ VGND VGND VPWR VPWR p_hh_pipe\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20006_ _01233_ VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__inv_2
XFILLER_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11710_ _02395_ _02524_ _02529_ VGND VGND VPWR VPWR _02648_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_87_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12690_ _03564_ _03615_ _03616_ _03614_ _03619_ VGND VGND VPWR VPWR _03620_ sky130_fd_sc_hd__o311a_1
X_11641_ net975 net692 net492 net698 VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__a22oi_4
XFILLER_70_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11572_ _02504_ net535 net658 net860 VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__a31o_1
X_14360_ _05262_ _05260_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__nand2_1
X_10523_ net1355 _01669_ _01670_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_118_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire701 a_h\[3\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__buf_6
X_13311_ net784 net986 net933 net787 VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__a22oi_2
XFILLER_11_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 a[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14291_ _01871_ net455 b_l\[14\] net709 _05193_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__o2111ai_4
X_10454_ _01617_ _01612_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__nand2_1
X_16030_ _06906_ _06895_ _06905_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__nand3_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13242_ net713 net923 net766 net710 VGND VGND VPWR VPWR _04157_ sky130_fd_sc_hd__and4_1
Xwire789 net792 VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__buf_12
Xwire778 net780 VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__buf_12
XFILLER_7_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10385_ term_mid\[33\] term_high\[33\] _01557_ _01482_ _01554_ VGND VGND VPWR VPWR
+ _01560_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_131_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13173_ _04087_ _04094_ _04095_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__a21oi_1
X_12124_ _03055_ net489 net687 VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__nand3_1
X_17981_ net627 net774 net769 net632 VGND VGND VPWR VPWR _08832_ sky130_fd_sc_hd__a22oi_1
XFILLER_69_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19720_ _00918_ _00922_ _00925_ _00921_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__o211ai_4
X_12055_ _02707_ _02862_ _02866_ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__o21ai_1
X_16932_ _07797_ _07798_ VGND VGND VPWR VPWR _07802_ sky130_fd_sc_hd__nand2_1
XFILLER_78_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11006_ _01947_ _01949_ _01944_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__a21o_1
X_16863_ net1103 _07694_ _07629_ _07627_ _07626_ VGND VGND VPWR VPWR _07733_ sky130_fd_sc_hd__a32oi_4
X_19651_ _00848_ _00851_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__nand2_2
X_15814_ net613 net521 VGND VGND VPWR VPWR _06693_ sky130_fd_sc_hd__nand2_1
X_18602_ net459 _07234_ _09369_ VGND VGND VPWR VPWR _09476_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_5_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19582_ _00776_ _00772_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__nor2_1
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16794_ _07537_ _07630_ _07659_ _07661_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__o22ai_2
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18533_ _09396_ _09387_ _09326_ _09398_ VGND VGND VPWR VPWR _09401_ sky130_fd_sc_hd__o211a_1
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15745_ _06586_ _06618_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__nand2_1
X_12957_ _03881_ _03882_ net665 net474 VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__nand4_1
XFILLER_45_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11908_ _02832_ _02839_ _02840_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__and3_1
X_15676_ _06507_ _06509_ _06553_ _06555_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__a22o_1
X_18464_ _09266_ _09291_ VGND VGND VPWR VPWR _09325_ sky130_fd_sc_hd__nand2_1
X_12888_ _03812_ _03813_ _09471_ _09668_ VGND VGND VPWR VPWR _03816_ sky130_fd_sc_hd__o2bb2a_1
X_11839_ _02773_ _02775_ net698 net1032 VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__nand4_1
X_17415_ _08277_ _08278_ _08273_ _08271_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__a31o_1
X_18395_ net769 net599 net593 net1123 VGND VGND VPWR VPWR _09250_ sky130_fd_sc_hd__a22o_1
X_14627_ _05384_ _05525_ _05524_ _05523_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__o211a_1
X_17346_ _08211_ _08206_ VGND VGND VPWR VPWR _08213_ sky130_fd_sc_hd__nand2_1
XFILLER_61_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14558_ _05435_ _05436_ _05455_ _05457_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__o22ai_2
X_17277_ _08000_ _08031_ _08140_ _08142_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__o22ai_4
X_13509_ _09155_ _09449_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__nor2_1
X_14489_ _05377_ _05378_ _05389_ _05390_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_134_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16228_ net570 net540 _07099_ _07102_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__a22oi_4
X_19016_ net592 net748 VGND VGND VPWR VPWR _09907_ sky130_fd_sc_hd__and2_1
X_16159_ _06912_ net1107 _07031_ net380 VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__a211oi_4
XTAP_TAPCELL_ROW_58_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19918_ _01120_ _01124_ _01132_ _01133_ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_95_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19849_ _01054_ _01056_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__nand3_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20624_ clknet_leaf_47_clk _00264_ VGND VGND VPWR VPWR p_ll_pipe\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_22_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20555_ clknet_leaf_18_clk _00195_ VGND VGND VPWR VPWR mid_sum\[18\] sky130_fd_sc_hd__dfxtp_1
X_20486_ clknet_leaf_45_clk _00126_ VGND VGND VPWR VPWR term_mid\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13860_ _04757_ _04760_ _04729_ _04759_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__o211ai_4
X_12811_ _09460_ _09668_ _03736_ _03737_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__o22a_1
X_13791_ _04581_ _04583_ _04694_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__a21o_1
XFILLER_103_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15530_ net627 net631 net532 net528 VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__nand4_2
X_12742_ net634 net514 net509 net638 VGND VGND VPWR VPWR _03672_ sky130_fd_sc_hd__a22o_1
X_12673_ _03244_ _03248_ _03115_ _03114_ _03247_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15461_ _06351_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__inv_2
X_11624_ _02435_ _02437_ _02560_ _02562_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__a2bb2oi_1
X_17200_ _08060_ _08065_ _08063_ VGND VGND VPWR VPWR _08068_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14412_ _09460_ _09471_ _04260_ _05133_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__o31a_1
X_18180_ net623 net759 VGND VGND VPWR VPWR _09027_ sky130_fd_sc_hd__nand2_1
X_15392_ _06238_ _06278_ _06284_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_41_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17131_ _07995_ _07996_ _07897_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__a21oi_4
X_11555_ _02361_ _02493_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__nand2_1
Xwire520 net524 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__buf_12
X_14343_ _05239_ _05241_ _05245_ _05116_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__o211ai_2
X_10506_ _01653_ _01657_ term_high\[55\] VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__and3_2
X_11486_ _02351_ _02353_ _02423_ _02424_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__o211ai_1
X_17062_ _09286_ _09613_ _07781_ _07925_ _07924_ VGND VGND VPWR VPWR _07931_ sky130_fd_sc_hd__o221ai_2
Xwire553 net555 VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__buf_12
XFILLER_11_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14274_ _05172_ _05145_ _05173_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__nand3_4
X_10437_ term_mid\[40\] term_high\[40\] term_mid\[41\] term_high\[41\] VGND VGND VPWR
+ VPWR _01604_ sky130_fd_sc_hd__a22o_1
X_16013_ _06889_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__inv_2
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13225_ net713 net710 _04133_ _04141_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__a31oi_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10368_ term_mid\[32\] term_high\[32\] VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__xor2_2
X_13156_ net265 _04075_ _04076_ _04077_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a2bb2oi_1
X_12107_ _03040_ _03041_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand2_1
X_17964_ net459 _06402_ _08815_ _08816_ VGND VGND VPWR VPWR _08817_ sky130_fd_sc_hd__o211a_1
XFILLER_69_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13087_ _04008_ _04009_ _04010_ _03970_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__a22o_1
X_10299_ term_low\[22\] term_mid\[22\] VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__nor2_1
XFILLER_111_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12038_ _02883_ _02888_ _02885_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a21oi_1
X_16915_ net578 net571 net513 net506 VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__and4_1
X_19703_ _09231_ _09362_ _00901_ _00904_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__o22a_1
X_17895_ _09340_ _09679_ _08751_ _08752_ VGND VGND VPWR VPWR _08754_ sky130_fd_sc_hd__o22a_1
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19634_ _00780_ _00828_ _00732_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_144_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16846_ _07703_ _07704_ _07712_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_0_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16777_ _07644_ _07647_ _07639_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19565_ net445 _00743_ _00745_ _00739_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__o31a_1
XFILLER_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13989_ net783 net650 net643 net788 VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__a22oi_1
XFILLER_34_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15728_ _06604_ _06607_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18516_ _09379_ _09372_ _09368_ _09378_ VGND VGND VPWR VPWR _09382_ sky130_fd_sc_hd__o211ai_2
X_19496_ _00631_ _00634_ _00681_ net1003 VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__a22oi_4
X_18447_ _09304_ _09306_ _09187_ _09189_ VGND VGND VPWR VPWR _09307_ sky130_fd_sc_hd__o2bb2ai_1
X_15659_ net542 net602 net624 net522 VGND VGND VPWR VPWR _06540_ sky130_fd_sc_hd__nand4_4
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18378_ _09151_ _09154_ _09149_ VGND VGND VPWR VPWR _09232_ sky130_fd_sc_hd__a21o_1
XFILLER_147_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17329_ net342 _08101_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__nand2_1
X_20340_ net793 net4 VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20271_ _01479_ _01510_ _01511_ _01515_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__o31a_1
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20607_ clknet_leaf_32_clk _00247_ VGND VGND VPWR VPWR p_ll_pipe\[5\] sky130_fd_sc_hd__dfxtp_1
X_11340_ net1062 _02278_ net671 net1024 _02277_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__o2111ai_4
X_20538_ clknet_leaf_38_clk net1364 VGND VGND VPWR VPWR mid_sum\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_116_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20469_ clknet_leaf_13_clk _00109_ VGND VGND VPWR VPWR term_high\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11271_ _02204_ _02207_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__nand2_1
XFILLER_118_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13010_ _03802_ _03803_ _03857_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__nand3_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10222_ net517 VGND VGND VPWR VPWR _09602_ sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_95_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16700_ _07442_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__nand2_1
XFILLER_48_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14961_ _05850_ _05853_ _05856_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__a21o_1
X_17680_ _08458_ _08462_ _08457_ VGND VGND VPWR VPWR _08544_ sky130_fd_sc_hd__o21ai_1
X_13912_ _04670_ net286 _04813_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__o21ai_1
X_14892_ _05789_ _05790_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16631_ _07393_ _07493_ _07500_ _07501_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__o211ai_1
XFILLER_114_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13843_ _04746_ _04748_ _04743_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__o21ai_2
X_16562_ _07297_ _07299_ _07298_ _07433_ _07432_ VGND VGND VPWR VPWR _07435_ sky130_fd_sc_hd__a32o_1
XFILLER_90_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19350_ _00524_ _00525_ _00526_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__a21o_1
X_10986_ _01927_ _01928_ _01914_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__a21o_1
X_18301_ net791 net582 VGND VGND VPWR VPWR _09148_ sky130_fd_sc_hd__nand2_1
X_13774_ _04586_ _04656_ _04658_ _04677_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__a31oi_4
X_15513_ _06398_ _06400_ net65 VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__a21oi_1
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16493_ _07263_ _07267_ _07363_ _07364_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__nand4_1
X_12725_ _03652_ _03653_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__nand2_1
X_19281_ _10043_ _10041_ _10045_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__o21a_4
XFILLER_31_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12656_ _03585_ _03586_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__nand2_1
X_18232_ _09053_ _09056_ _09075_ VGND VGND VPWR VPWR _09079_ sky130_fd_sc_hd__o21ai_2
XFILLER_70_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15444_ _06301_ _06306_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__o21ai_1
XFILLER_128_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11607_ _02541_ _02542_ _02478_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__nand3_2
X_18163_ _09005_ _08954_ _09004_ VGND VGND VPWR VPWR _09011_ sky130_fd_sc_hd__nand3_1
X_12587_ _09504_ _03510_ _03421_ _03512_ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__o211a_1
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15375_ _06265_ _06266_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__nand2_1
XFILLER_129_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17114_ _07980_ _07981_ _07978_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__o21ai_4
X_14326_ _05050_ _05065_ _05225_ _05063_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__o211a_1
XFILLER_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11538_ _02390_ _02416_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__nand2_1
X_18094_ _08940_ _08942_ VGND VGND VPWR VPWR _08943_ sky130_fd_sc_hd__nand2_1
Xhold408 p_ll\[20\] VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _02254_ _02257_ _02258_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__a21boi_2
XFILLER_116_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17045_ _07906_ _07908_ _07913_ _07815_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__a22oi_1
Xhold419 p_ll_pipe\[18\] VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_14257_ _04988_ _05159_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__nand2_2
X_13208_ _04126_ _04123_ net198 VGND VGND VPWR VPWR _04129_ sky130_fd_sc_hd__a21oi_1
X_14188_ _05084_ _05086_ _05091_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__a21o_1
XFILLER_124_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13139_ _04017_ _04060_ _04062_ _04059_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__a22o_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ net609 net732 VGND VGND VPWR VPWR _09887_ sky130_fd_sc_hd__nand2_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17947_ _08770_ _08791_ VGND VGND VPWR VPWR _08804_ sky130_fd_sc_hd__nor2_1
Xclone251 net674 VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__clkbuf_16
X_17878_ _09297_ _09679_ _08692_ _08693_ VGND VGND VPWR VPWR _08738_ sky130_fd_sc_hd__o31a_1
X_16829_ _07698_ _07628_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__nand2_1
Xclone273 net528 net532 VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__nand2_4
Xclone262 net524 VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__clkbuf_16
X_19617_ _00812_ _00793_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__nand2_1
XFILLER_38_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19548_ _09264_ _09297_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__nor2_1
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19479_ _00661_ _00662_ _00664_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__a21o_1
XFILLER_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20323_ net793 net20 VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__and2_1
XFILLER_143_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap672 net674 VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__buf_12
Xmax_cap650 net870 VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__buf_12
X_20254_ _01350_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__nand2_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap661 a_h\[10\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__buf_12
XFILLER_135_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap683 net932 VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__buf_8
Xmax_cap694 net695 VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__buf_6
XFILLER_0_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20185_ _01423_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__and2b_1
XFILLER_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10840_ net795 net1157 VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__and2_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10771_ _01787_ _01789_ _01796_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__a21oi_1
XFILLER_53_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12510_ _09482_ _09613_ _03128_ _03261_ VGND VGND VPWR VPWR _03442_ sky130_fd_sc_hd__o22a_1
X_13490_ _04353_ _04357_ _04358_ _04345_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_9_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12441_ _03373_ _03123_ _03247_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_97_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12372_ _03302_ _03303_ _09417_ _09668_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15160_ _05994_ _05995_ _06050_ _06051_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__a22o_1
XFILLER_126_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11323_ _02261_ _02262_ _02252_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__nand3_2
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15091_ _05902_ _05968_ _05969_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__a21o_1
X_14111_ _05013_ _05014_ _05010_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__a21o_1
X_11254_ net702 net697 net1018 net507 _02189_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__a41o_1
X_14042_ _04940_ _04946_ _04945_ _04869_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__o211ai_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18850_ _09692_ _09694_ _09688_ VGND VGND VPWR VPWR _09742_ sky130_fd_sc_hd__a21boi_2
X_10205_ net696 VGND VGND VPWR VPWR _09417_ sky130_fd_sc_hd__inv_8
X_11185_ _02122_ _02124_ _02123_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_128_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17801_ _08661_ _08659_ _08657_ VGND VGND VPWR VPWR _08663_ sky130_fd_sc_hd__nand3_1
XFILLER_121_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15993_ _09275_ _09581_ net1070 _06867_ _06865_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__o221ai_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18781_ _09651_ _09667_ _09669_ VGND VGND VPWR VPWR _09672_ sky130_fd_sc_hd__nand3_1
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17732_ _08515_ _08512_ _08510_ _08507_ VGND VGND VPWR VPWR _08595_ sky130_fd_sc_hd__o2bb2ai_1
X_14944_ _09449_ _09460_ net455 _05835_ _05837_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_141_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17663_ _08524_ _08526_ _08478_ VGND VGND VPWR VPWR _08527_ sky130_fd_sc_hd__a21o_1
X_16614_ _07483_ _07484_ _07485_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__a21o_1
XFILLER_63_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14875_ _05771_ _05774_ _05773_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nand3b_4
X_19402_ _00583_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__inv_2
XFILLER_36_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17594_ _08270_ _08367_ _08365_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__a21o_1
XFILLER_63_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13826_ net1122 net667 VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__nand2_1
X_16545_ _07342_ _07343_ _07415_ _07416_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__a22o_1
X_10969_ _01885_ _01890_ _01889_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__o21ai_4
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13757_ _09177_ _09308_ _01860_ _04555_ _04663_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__o221a_1
X_19333_ net603 net729 net725 net609 VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__a22o_1
X_16476_ _07256_ _07279_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__nand2_1
X_12708_ net648 net500 VGND VGND VPWR VPWR _03638_ sky130_fd_sc_hd__nand2_1
X_19264_ net765 net562 VGND VGND VPWR VPWR _10165_ sky130_fd_sc_hd__nand2_1
XFILLER_31_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18215_ net782 net585 VGND VGND VPWR VPWR _09062_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_61_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ _04593_ _04594_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__nand2_2
X_15427_ _06274_ _06318_ _06271_ _06272_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__and4_1
X_12639_ _03532_ _03533_ _03568_ _03569_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_61_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19195_ _10087_ _10088_ VGND VGND VPWR VPWR _10091_ sky130_fd_sc_hd__nand2_2
XFILLER_129_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18146_ _08990_ _08988_ _08989_ VGND VGND VPWR VPWR _08994_ sky130_fd_sc_hd__a21oi_2
X_15358_ _06189_ _06196_ _06197_ _06190_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__a31o_4
X_18077_ _09155_ _09199_ net459 _06681_ _08920_ VGND VGND VPWR VPWR _08926_ sky130_fd_sc_hd__o221ai_4
X_14309_ _05057_ _05200_ _05209_ _05210_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__o211ai_4
X_15289_ _06101_ _06105_ _06113_ _06104_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17028_ _07777_ _07843_ _07841_ _07834_ VGND VGND VPWR VPWR _07897_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18979_ _09771_ _09845_ _09844_ VGND VGND VPWR VPWR _09870_ sky130_fd_sc_hd__a21boi_4
XFILLER_39_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer313 _06593_ VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__buf_1
Xrebuffer302 net1095 VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer324 b_l\[6\] VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer335 _04737_ VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20306_ _01540_ _01549_ _01551_ _01502_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__o22ai_1
XPHY_EDGE_ROW_141_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap480 b_h\[13\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__buf_8
Xmax_cap491 net492 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_6
XFILLER_89_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20237_ _01437_ _01477_ _01479_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__nand3_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20168_ _09286_ _09384_ _01385_ _01388_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__o31ai_1
XFILLER_130_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12990_ _03914_ _03916_ _03900_ VGND VGND VPWR VPWR _03917_ sky130_fd_sc_hd__nand3_1
X_20099_ _01324_ _01331_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_123_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ net358 _02873_ _02874_ _02708_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a211o_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11872_ _02805_ _02806_ _02693_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__nand3_2
X_14660_ _05286_ _05452_ net427 _05559_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10823_ _01839_ _01840_ _01841_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__a21oi_1
X_13611_ net785 net666 net660 net1058 VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__a22oi_4
X_14591_ _05313_ _05314_ _05311_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__a21oi_1
X_16330_ _02588_ net848 _07203_ VGND VGND VPWR VPWR _07204_ sky130_fd_sc_hd__a21oi_1
X_13542_ _04451_ net352 _04438_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__a21o_1
XFILLER_53_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10754_ p_hl\[19\] p_lh\[19\] _01767_ _01781_ _01780_ VGND VGND VPWR VPWR _01782_
+ sky130_fd_sc_hd__a221o_1
X_16261_ _09199_ _09613_ _07134_ _07135_ VGND VGND VPWR VPWR _07136_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_101_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18000_ _08826_ _08848_ _08849_ _08850_ VGND VGND VPWR VPWR _08851_ sky130_fd_sc_hd__and4_1
X_13473_ _04314_ _04317_ _04383_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__nand3_1
X_10685_ p_hl\[10\] p_lh\[10\] VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__nor2_1
X_16192_ net620 net496 net491 net841 VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__a22oi_4
X_12424_ _03252_ _03355_ _03356_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__nand3b_4
X_15212_ net1025 net657 _05043_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__and3_1
XFILLER_138_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12355_ _02998_ _03157_ net985 _03284_ VGND VGND VPWR VPWR _03288_ sky130_fd_sc_hd__o2bb2ai_4
X_15143_ _06039_ _05912_ _06038_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_134_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11306_ net361 _02205_ _02242_ _02243_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__a211o_1
XFILLER_5_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12286_ _03218_ _03219_ VGND VGND VPWR VPWR _03220_ sky130_fd_sc_hd__nand2_1
X_19951_ _01166_ _01168_ _01170_ VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__and3_1
X_15074_ _05970_ _05902_ _05968_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__nand3_1
X_11237_ _02177_ net362 VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__nand2_1
X_18902_ _09789_ _09790_ VGND VGND VPWR VPWR _09794_ sky130_fd_sc_hd__nand2_1
X_19882_ net895 net549 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__nand2_1
X_14025_ _04927_ net689 net746 VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__nand3_1
X_11168_ net707 net702 net1018 net507 _02109_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__a41o_1
X_18833_ _09574_ _09723_ _09719_ VGND VGND VPWR VPWR _09726_ sky130_fd_sc_hd__a21oi_2
X_18764_ _09484_ _09487_ VGND VGND VPWR VPWR _09653_ sky130_fd_sc_hd__nand2_1
X_15976_ _06850_ _06852_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__nor2_1
X_11099_ _02042_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__inv_2
X_17715_ _08575_ _08576_ _08561_ VGND VGND VPWR VPWR _08578_ sky130_fd_sc_hd__a21o_1
X_18695_ _09414_ _09415_ net185 _09573_ _09572_ VGND VGND VPWR VPWR _09578_ sky130_fd_sc_hd__o221ai_4
X_14927_ net730 net668 VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__nand2_1
X_17646_ _08509_ _08380_ VGND VGND VPWR VPWR _08510_ sky130_fd_sc_hd__nand2_1
X_14858_ net285 _05633_ _05753_ net1011 net715 VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__a32o_1
XFILLER_35_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_91_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17577_ _08438_ _08440_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_63_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13809_ _04635_ net683 net757 VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__nand3_1
X_16528_ net307 _07389_ _07399_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__a21o_1
X_19316_ _00488_ _00490_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__nand2_1
X_14789_ _05683_ _05685_ _05680_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__a21o_1
XFILLER_32_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16459_ _07194_ _07198_ _07328_ _07329_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__a22oi_2
X_19247_ _10142_ _10144_ VGND VGND VPWR VPWR _10147_ sky130_fd_sc_hd__nand2_1
X_19178_ net369 _09890_ _09893_ VGND VGND VPWR VPWR _10073_ sky130_fd_sc_hd__a21oi_1
XFILLER_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18129_ _08916_ _08921_ VGND VGND VPWR VPWR _08977_ sky130_fd_sc_hd__nand2_1
XFILLER_117_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20022_ _01202_ _01249_ _01250_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__nand3_2
XFILLER_101_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer20 b_l\[1\] VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_27_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer31 b_h\[10\] VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer42 net1039 VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_15_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer64 a_h\[8\] VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__clkbuf_2
Xrebuffer53 _10058_ VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__clkbuf_2
Xrebuffer75 net654 VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer97 net893 VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__buf_4
Xrebuffer86 b_l\[2\] VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20786_ clknet_leaf_25_clk _00426_ VGND VGND VPWR VPWR a_l\[8\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_12_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10470_ term_mid\[46\] term_high\[46\] _01631_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__a21o_1
XFILLER_136_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer132 a_l\[5\] VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer110 a_h\[13\] VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__buf_2
Xrebuffer121 b_l\[10\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer154 _02677_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer143 a_l\[15\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer165 net960 VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__buf_1
Xrebuffer176 net972 VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12140_ _03070_ _03072_ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__nor2_1
XFILLER_108_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer187 _00467_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd1_1
X_12071_ net906 net518 VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__nand2_1
Xhold580 p_lh\[31\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11022_ _09417_ _09592_ _01919_ _01962_ _01961_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__o221ai_2
X_15830_ _06674_ _06705_ _06706_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__nand3_4
XFILLER_66_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15761_ _06634_ _06636_ _06508_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__nand3_2
X_12973_ _03896_ _03898_ VGND VGND VPWR VPWR _03900_ sky130_fd_sc_hd__nor2_1
X_11924_ _02752_ _02859_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__nand2_1
X_15692_ _06504_ _06572_ _06571_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__a21oi_1
X_17500_ _08362_ _08363_ _08364_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__a21o_1
X_18480_ _09333_ _09336_ _09327_ _09338_ VGND VGND VPWR VPWR _09343_ sky130_fd_sc_hd__o211ai_2
XFILLER_45_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14712_ net736 net670 VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_103_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _08295_ _08221_ _08227_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__nor3_1
X_14643_ _05468_ _05471_ _05495_ _05542_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__o211ai_1
X_11855_ _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__inv_2
XFILLER_72_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11786_ net653 net526 net1059 net658 VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__a22oi_1
X_10806_ p_hl\[27\] p_lh\[27\] VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__xor2_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17362_ _08221_ _08227_ _08226_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__o21ai_2
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19101_ _09976_ _09977_ _09984_ _09986_ VGND VGND VPWR VPWR _09992_ sky130_fd_sc_hd__nand4_1
X_14574_ _05472_ _05474_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_31_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16313_ _07088_ _07156_ _07154_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__a21oi_1
X_17293_ _08020_ _08030_ _08160_ VGND VGND VPWR VPWR _08161_ sky130_fd_sc_hd__a21oi_1
X_10737_ _01765_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__nor2_1
X_13525_ _04430_ _04431_ _04399_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_136_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16244_ _07112_ _07117_ _07115_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__a21oi_2
X_13456_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__nand2_1
X_19032_ _09920_ net1101 _09917_ VGND VGND VPWR VPWR _09923_ sky130_fd_sc_hd__nand3b_2
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12407_ _03339_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__inv_2
X_10668_ p_hl\[7\] p_lh\[7\] VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__nand2_1
XFILLER_9_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 net107 VGND VGND VPWR VPWR p[47] sky130_fd_sc_hd__buf_2
X_16175_ _06950_ _07047_ net154 VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__nand3_4
X_10599_ _09690_ net1227 VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__and2_1
X_13387_ _04278_ _04279_ _04295_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__o21ai_1
Xoutput118 net118 VGND VGND VPWR VPWR p[57] sky130_fd_sc_hd__buf_2
Xoutput129 net129 VGND VGND VPWR VPWR p[9] sky130_fd_sc_hd__buf_2
X_12338_ _03256_ _03266_ _03267_ _03269_ _03253_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__a32o_1
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15126_ _06019_ _06020_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__nand2_2
XFILLER_142_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12269_ _03045_ _03046_ _03060_ _03062_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__o31a_1
X_19934_ _01000_ _01047_ _01153_ _01154_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__nand4_4
X_15057_ _05922_ _05951_ _05952_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_56_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14008_ _04888_ _04907_ _04873_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__a21oi_1
X_19865_ _00858_ _00965_ _00966_ _00979_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__a31oi_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18816_ _09707_ _09708_ VGND VGND VPWR VPWR _09709_ sky130_fd_sc_hd__nand2_1
X_19796_ _01005_ _01006_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15959_ net173 _06836_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__nand2_1
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18747_ _09632_ _09633_ VGND VGND VPWR VPWR _09634_ sky130_fd_sc_hd__nand2_2
XFILLER_49_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18678_ _09412_ _09553_ _09555_ VGND VGND VPWR VPWR _09560_ sky130_fd_sc_hd__and3_1
XFILLER_36_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17629_ _08490_ _08491_ VGND VGND VPWR VPWR _08493_ sky130_fd_sc_hd__nand2_1
X_20640_ clknet_leaf_18_clk _00280_ VGND VGND VPWR VPWR p_hh\[6\] sky130_fd_sc_hd__dfxtp_1
X_20571_ clknet_leaf_26_clk _00211_ VGND VGND VPWR VPWR p_hh_pipe\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20005_ _01228_ _01229_ _01230_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__nand3_4
XFILLER_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11640_ net706 net487 VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__nand2_2
X_11571_ _02509_ _02500_ _02495_ _02508_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__o211ai_2
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10522_ net1355 _01669_ net65 VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__a21oi_1
X_13310_ net787 net784 net986 net933 VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nand4_4
Xwire724 net1095 VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__buf_6
X_20769_ clknet_leaf_59_clk _00409_ VGND VGND VPWR VPWR a_h\[7\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_118_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14290_ _05193_ net709 b_l\[14\] _05192_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__and4_2
X_10453_ _01595_ _01616_ _01615_ _01612_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__a211o_1
XFILLER_136_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13241_ _09690_ _04155_ _04156_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__and3_1
X_10384_ _01417_ _01460_ _01513_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__a31o_1
XFILLER_123_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13172_ _04087_ _04094_ net793 VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_131_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12123_ _03053_ _03055_ _09428_ _09646_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__o2bb2ai_1
X_17980_ net774 net769 _06401_ VGND VGND VPWR VPWR _08831_ sky130_fd_sc_hd__and3_1
X_12054_ _02707_ _02862_ _02866_ VGND VGND VPWR VPWR _02989_ sky130_fd_sc_hd__o21a_1
X_16931_ _07790_ _07796_ _07798_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__a21oi_2
XFILLER_78_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11005_ _01944_ _01947_ _01949_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__nand3_1
X_16862_ _07587_ _07731_ _07732_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__o21ba_1
X_19650_ _00845_ _00847_ _00850_ _00702_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__a22oi_1
X_15813_ net1127 net515 VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__nand2_2
X_16793_ _07662_ _07631_ _07660_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__nand3_4
X_18601_ _09365_ _09380_ _09382_ VGND VGND VPWR VPWR _09475_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_5_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19581_ _00770_ _00771_ _00774_ _00646_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__o2bb2ai_4
X_15744_ _06585_ _06622_ _06621_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__nand3_4
X_18532_ net303 _09347_ _09386_ _09393_ VGND VGND VPWR VPWR _09400_ sky130_fd_sc_hd__o211ai_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12956_ _03881_ _03882_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__nand2_1
X_11907_ _02832_ _02841_ _02842_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__nand3b_4
X_15675_ _06549_ _06552_ _06510_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__o21bai_2
X_18463_ _09290_ _09295_ net252 _09296_ VGND VGND VPWR VPWR _09324_ sky130_fd_sc_hd__a2bb2oi_2
X_12887_ _02362_ _02589_ net944 net478 _03812_ VGND VGND VPWR VPWR _03815_ sky130_fd_sc_hd__o2111ai_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11838_ net692 net687 net497 net492 VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__nand4_2
X_17414_ _08269_ _08270_ _08280_ VGND VGND VPWR VPWR _08281_ sky130_fd_sc_hd__a21o_1
X_18394_ net1146 net599 net593 net1123 VGND VGND VPWR VPWR _09249_ sky130_fd_sc_hd__a22oi_1
X_14626_ _05523_ _05524_ _05526_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__a21o_1
X_17345_ _09319_ _09613_ _08052_ _08210_ _08208_ VGND VGND VPWR VPWR _08212_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_44_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _05437_ _05456_ _05458_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__nand3_1
XFILLER_20_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11769_ _02649_ _02705_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_40_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_8
X_13508_ _04412_ _04413_ _04416_ _04349_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_146_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17276_ _08000_ _08031_ _08141_ _08143_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__a2bb2oi_1
X_19015_ _09904_ _09905_ VGND VGND VPWR VPWR _09906_ sky130_fd_sc_hd__nand2_2
X_14488_ _05385_ _05386_ _05388_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__a21oi_1
XFILLER_146_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16227_ net582 net572 net532 net528 VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__nand4_4
XTAP_TAPCELL_ROW_58_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13439_ net785 net675 net673 net1058 VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__a22oi_4
X_16158_ net1107 _06912_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15109_ _06005_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__inv_2
XFILLER_142_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16089_ _09188_ _09613_ _06898_ _06961_ _06960_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_71_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19917_ _01134_ _01124_ net332 VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__nand3_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19848_ _01061_ _01062_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__nand2_2
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19779_ _00871_ _00876_ _00875_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_69_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20623_ clknet_leaf_47_clk _00263_ VGND VGND VPWR VPWR p_ll_pipe\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_31_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20554_ clknet_leaf_18_clk _00194_ VGND VGND VPWR VPWR mid_sum\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20485_ clknet_leaf_44_clk _00125_ VGND VGND VPWR VPWR term_mid\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12810_ _02278_ _02589_ net674 net478 _03738_ VGND VGND VPWR VPWR _03739_ sky130_fd_sc_hd__o2111a_2
XTAP_TAPCELL_ROW_2_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13790_ _04581_ _04583_ _04697_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__and3_1
X_12741_ _03430_ _03507_ _03511_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__o21ai_1
X_12672_ _03372_ _03496_ VGND VGND VPWR VPWR _03603_ sky130_fd_sc_hd__nor2_2
X_15460_ _06315_ _06349_ net388 VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__nand3_1
X_11623_ _02431_ _02445_ _02558_ _02559_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__o211ai_2
X_14411_ net746 _05125_ net676 _05127_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__a31o_1
X_17130_ _07989_ _07991_ _07996_ _07897_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__o211ai_1
Xclkbuf_leaf_22_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_15391_ _06282_ net657 net716 VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_41_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11554_ _02357_ _02364_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__nand2_1
X_14342_ _05242_ _05245_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nand2_1
X_10505_ _01653_ _01657_ net1347 VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__a21oi_1
X_11485_ _02423_ _02424_ net269 VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__a21bo_1
X_17061_ _07924_ _07927_ _07921_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__a21o_1
X_14273_ _05169_ net314 _05146_ _05175_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__o211ai_4
X_10436_ term_mid\[42\] term_high\[42\] VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__xor2_1
X_16012_ _06883_ _06884_ _06874_ _06875_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__o211ai_4
X_13224_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__nor2_1
XFILLER_124_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13155_ net266 _04075_ _04076_ _04077_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__and4bb_1
X_10367_ _01375_ _01386_ _01397_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__o21a_1
X_12106_ net692 net483 VGND VGND VPWR VPWR _03041_ sky130_fd_sc_hd__nand2_1
X_17963_ _08813_ _08814_ net779 net632 VGND VGND VPWR VPWR _08816_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_53_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _03968_ _03969_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__o21ai_1
X_10298_ net794 _00644_ _00655_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__and3_1
X_12037_ _02886_ _02890_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__nand2_1
X_16914_ net571 net506 VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__nand2_1
XFILLER_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19702_ _00905_ net718 net598 _00903_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__and4_2
X_17894_ _09340_ _09679_ _08751_ _08752_ VGND VGND VPWR VPWR _08753_ sky130_fd_sc_hd__nor4_1
X_19633_ _00777_ _00779_ _00828_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_144_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16845_ _07704_ _07712_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16776_ net558 net874 net534 net530 VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__nand4_4
XFILLER_81_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19564_ _00755_ net445 _00740_ _00753_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__o211ai_2
XFILLER_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13988_ net783 net650 VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__nand2_1
X_15727_ a_l\[4\] net607 net531 net527 VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__nand4_2
X_12939_ _03862_ _03866_ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__and2_1
X_18515_ _09379_ _09372_ _09367_ _09378_ VGND VGND VPWR VPWR _09381_ sky130_fd_sc_hd__o211ai_1
XFILLER_61_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19495_ _00681_ _00634_ _00631_ _00682_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__nand4_4
X_15658_ _06536_ _06537_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__nand2_1
X_18446_ _09302_ _09215_ _09301_ VGND VGND VPWR VPWR _09306_ sky130_fd_sc_hd__nand3_4
X_14609_ _05334_ net390 _05362_ _05369_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__and4_1
XFILLER_33_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
X_15589_ _09166_ _09602_ _06466_ _06469_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__o211ai_2
X_18377_ _09162_ _09228_ VGND VGND VPWR VPWR _09230_ sky130_fd_sc_hd__nand2_1
XFILLER_146_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17328_ _08187_ _08189_ _08191_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__nand3_2
XFILLER_146_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17259_ _07965_ _08089_ _08123_ _08124_ VGND VGND VPWR VPWR _08127_ sky130_fd_sc_hd__o211a_1
XFILLER_108_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20270_ _01512_ _01514_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__a21oi_1
XFILLER_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_110_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20606_ clknet_leaf_32_clk _00246_ VGND VGND VPWR VPWR p_ll_pipe\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20537_ clknet_leaf_38_clk net1327 VGND VGND VPWR VPWR mid_sum\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20468_ clknet_leaf_14_clk _00108_ VGND VGND VPWR VPWR term_high\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_134_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11270_ _02209_ _02211_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__nand2_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10221_ net536 VGND VGND VPWR VPWR _09592_ sky130_fd_sc_hd__clkinv_8
XPHY_EDGE_ROW_18_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20399_ clknet_leaf_46_clk _00039_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14960_ _05850_ _05853_ _05856_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__nand3_1
XFILLER_102_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13911_ _04815_ _04812_ net164 VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__o21ai_1
X_14891_ _09384_ _09428_ _05785_ _05787_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_126_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ _07395_ _07500_ _07501_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__nand3_2
XFILLER_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13842_ net788 net783 net656 net650 VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__nand4_2
X_16561_ _07302_ _07432_ _07433_ VGND VGND VPWR VPWR _07434_ sky130_fd_sc_hd__nand3_2
XFILLER_74_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13773_ _04487_ _04550_ _04584_ _04678_ _04679_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__o2111ai_4
XFILLER_16_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10985_ _01927_ _01928_ _01914_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__nand3_1
X_18300_ _09068_ _09072_ VGND VGND VPWR VPWR _09147_ sky130_fd_sc_hd__nand2_1
XFILLER_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12724_ _03653_ VGND VGND VPWR VPWR _03654_ sky130_fd_sc_hd__inv_2
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19280_ _10041_ _10043_ _10045_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__o21ai_2
X_15512_ _06369_ _06370_ _06387_ _06389_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__o22a_1
X_16492_ _07363_ _07364_ _07352_ VGND VGND VPWR VPWR _07365_ sky130_fd_sc_hd__a21o_1
X_18231_ net372 _09073_ _09074_ _09057_ VGND VGND VPWR VPWR _09078_ sky130_fd_sc_hd__o211ai_4
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12655_ _09428_ _09679_ _03582_ _03583_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__o211ai_4
X_15443_ net162 VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__inv_2
X_11606_ _02543_ _02544_ _02479_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__a21oi_4
XFILLER_90_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18162_ _08954_ _09005_ VGND VGND VPWR VPWR _09010_ sky130_fd_sc_hd__nand2_2
X_12586_ _03516_ VGND VGND VPWR VPWR _03517_ sky130_fd_sc_hd__inv_2
X_15374_ net726 net722 net642 net640 VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__nand4_1
X_11537_ _02471_ _02472_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__nand2_1
X_17113_ _07976_ _07977_ _07948_ VGND VGND VPWR VPWR _07982_ sky130_fd_sc_hd__a21o_1
X_18093_ _08935_ _08938_ _08899_ VGND VGND VPWR VPWR _08942_ sky130_fd_sc_hd__nand3_1
X_14325_ _05223_ _05224_ _05227_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__nand3_1
Xwire351 _04755_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_1
XFILLER_144_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_139_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17044_ _07819_ _07822_ _07652_ _07816_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__o22ai_4
Xhold409 term_low\[10\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11468_ _02294_ net439 _02402_ _02405_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o211ai_2
X_14256_ net783 net639 net636 net788 VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_36_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10419_ term_mid\[40\] term_high\[40\] VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__nor2_1
X_11399_ net983 net706 net975 net492 VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__and4_1
XFILLER_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13207_ _04111_ _04122_ _04125_ _04094_ net198 VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__o221ai_1
X_14187_ _05084_ _05090_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__nand2_1
XFILLER_98_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13138_ _04022_ _04019_ _04058_ _04057_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a22o_1
X_18995_ net603 net598 net1091 net738 VGND VGND VPWR VPWR _09886_ sky130_fd_sc_hd__nand4_2
X_17946_ _08769_ _08788_ _08789_ VGND VGND VPWR VPWR _08803_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_2_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
X_13069_ _03990_ _03991_ _03992_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__nand3_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17877_ _08694_ _08732_ _08734_ _08698_ VGND VGND VPWR VPWR _08737_ sky130_fd_sc_hd__and4_1
X_16828_ _07624_ _07625_ _07697_ _07696_ VGND VGND VPWR VPWR _07699_ sky130_fd_sc_hd__o211ai_2
XFILLER_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclone252 net641 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__clkbuf_16
XFILLER_54_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19616_ _00790_ _00792_ _00808_ _00811_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__o211ai_2
XFILLER_80_102 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone296 a_l\[10\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__clkbuf_16
Xclone285 net1092 VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_45_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19547_ _10170_ _00637_ _00639_ _00636_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__a22o_1
X_16759_ _07522_ _07531_ _07532_ _07519_ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__a31oi_1
XTAP_TAPCELL_ROW_66_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19478_ _00661_ _00662_ _00664_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__a21oi_1
X_18429_ net457 _06480_ _09123_ _09282_ _09283_ VGND VGND VPWR VPWR _09288_ sky130_fd_sc_hd__o2111ai_4
XFILLER_22_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20322_ net793 net19 VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__and2_1
XFILLER_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap651 net868 VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__buf_6
Xmax_cap640 net912 VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__buf_8
X_20253_ _01351_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__and2_1
Xmax_cap662 net663 VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_110_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap684 a_h\[6\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__buf_12
Xmax_cap673 net674 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__clkbuf_8
Xmax_cap695 net1009 VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__buf_8
X_20184_ _01367_ net329 _01419_ _01420_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__nand4_1
XFILLER_130_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_103_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10770_ p_hl\[21\] p_lh\[21\] _01795_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_121_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12440_ _03112_ _03113_ _03244_ _03248_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_138_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12371_ _03303_ net475 net696 _03302_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__and4_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14110_ _05013_ _05014_ net746 net683 VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__nand4_2
X_11322_ _02253_ _02259_ _02260_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__nand3_2
XFILLER_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15090_ _05985_ _05986_ _05987_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__o21a_1
X_11253_ net708 net501 _02192_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__a22o_1
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14041_ _04768_ _04870_ _04941_ _04942_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__o211ai_4
XFILLER_106_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10204_ net700 VGND VGND VPWR VPWR _09406_ sky130_fd_sc_hd__inv_8
X_11184_ _02120_ _02121_ _02125_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_128_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17800_ _08520_ _08590_ _08605_ _08660_ VGND VGND VPWR VPWR _08662_ sky130_fd_sc_hd__o211ai_2
X_15992_ a_l\[7\] net1116 net531 net527 VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__nand4_1
X_18780_ _09647_ _09648_ _09670_ VGND VGND VPWR VPWR _09671_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17731_ net1072 net472 VGND VGND VPWR VPWR _08594_ sky130_fd_sc_hd__nand2_1
X_14943_ _05836_ _05838_ net720 net685 VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_141_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17662_ _08520_ _08522_ _08382_ _08424_ VGND VGND VPWR VPWR _08526_ sky130_fd_sc_hd__o2bb2ai_2
X_14874_ net163 _05655_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__nand2_1
XFILLER_36_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16613_ _07332_ _07320_ _07331_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__o21ai_2
X_13825_ _04730_ _04731_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__nand2_2
X_19401_ _00508_ _00511_ _00524_ _00581_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__o211ai_2
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_106_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17593_ _08456_ _08457_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__nand2_1
X_16544_ _07347_ _07416_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__nand2_1
X_10968_ net466 _01912_ _01913_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_106_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13756_ net741 net734 net709 net703 VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_48_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19332_ net887 net603 net729 net725 VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__nand4_1
X_16475_ _07342_ _07343_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__nand2_1
X_12707_ net872 b_h\[10\] VGND VGND VPWR VPWR _03637_ sky130_fd_sc_hd__nand2_1
X_19263_ _09816_ net549 net881 VGND VGND VPWR VPWR _10164_ sky130_fd_sc_hd__and3_1
X_13687_ net1064 net660 net656 net788 VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__a22oi_4
X_12638_ _03563_ _03565_ _03566_ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__nand3_2
X_18214_ net779 net1113 VGND VGND VPWR VPWR _09061_ sky130_fd_sc_hd__nand2_1
X_10899_ net794 net1337 VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__and2_1
X_15426_ _06265_ _06266_ _06269_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__o21ai_1
X_19194_ net592 net1092 net738 net598 VGND VGND VPWR VPWR _10090_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_139_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12569_ _03465_ _03470_ _03469_ VGND VGND VPWR VPWR _03500_ sky130_fd_sc_hd__a21bo_1
X_18145_ _08986_ _08988_ _08983_ VGND VGND VPWR VPWR _08993_ sky130_fd_sc_hd__a21oi_2
X_15357_ _06247_ _06248_ _06240_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__nand3_2
XFILLER_129_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18076_ _08920_ _08921_ _08916_ VGND VGND VPWR VPWR _08925_ sky130_fd_sc_hd__a21o_1
X_14308_ _05206_ _05208_ _05203_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__a21o_1
X_15288_ _06111_ _06112_ _06101_ _06105_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__o22a_1
X_17027_ _07834_ _07841_ _07843_ _07777_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__a2bb2oi_2
X_14239_ _05140_ _05142_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__nand2_1
XFILLER_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18978_ _09771_ _09845_ _09843_ _09840_ VGND VGND VPWR VPWR _09869_ sky130_fd_sc_hd__o2bb2ai_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17929_ _08779_ _08786_ VGND VGND VPWR VPWR _08787_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_53_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_135_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer336 _04461_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__buf_8
Xrebuffer325 net768 VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__buf_2
XFILLER_147_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20305_ _01522_ _01523_ _01539_ net158 VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__a211o_1
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap470 _01562_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_92_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap481 b_h\[13\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_8
XFILLER_103_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap492 net495 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_12
X_20236_ _01436_ _01434_ _01479_ _01477_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__a2bb2o_2
X_20167_ net794 _01405_ _01406_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__and3_1
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20098_ _01321_ _01323_ _01329_ _01330_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__nand4_1
X_11940_ net358 _02873_ _02875_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_123_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11871_ _02803_ net949 _02698_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a21oi_2
XFILLER_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10822_ _01839_ _01840_ net795 VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__o21ai_1
X_13610_ net789 net660 VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__nand2_1
X_14590_ _05312_ _05319_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__nand2_1
X_10753_ p_hl\[17\] p_lh\[17\] _01769_ _01774_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__o211a_1
XFILLER_71_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13541_ _04342_ _04446_ _04447_ _04449_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__nand4_4
XFILLER_13_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16260_ _06961_ net512 net966 VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_101_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13472_ _04381_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__nand2_1
X_10684_ _01721_ _01722_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__nor2_1
X_15211_ net726 net657 VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__nand2_1
X_16191_ net629 net487 VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__nand2_1
X_12423_ _03346_ _03347_ _03352_ _03353_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__nand4_1
X_12354_ _02899_ _02996_ _03157_ _03285_ VGND VGND VPWR VPWR _03287_ sky130_fd_sc_hd__o211ai_4
X_15142_ _06012_ _06014_ _06034_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_134_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ _02242_ _02243_ _02245_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__o21ai_1
X_19950_ _01160_ _01162_ _01086_ _01171_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__a31o_4
X_15073_ _05968_ _05970_ _05902_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__a21oi_2
X_12285_ _03124_ _03216_ _03217_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__nand3_4
X_18901_ _09791_ _09792_ VGND VGND VPWR VPWR _09793_ sky130_fd_sc_hd__nand2_1
X_14024_ _09264_ _09428_ _04708_ _04925_ _04924_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__o221ai_2
XFILLER_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11236_ _02176_ _02177_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__nand2_1
X_19881_ _00872_ _00982_ _00987_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__o21ai_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11167_ net712 net501 _02106_ _02108_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__a22o_1
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18832_ _09719_ _09721_ _09724_ VGND VGND VPWR VPWR _09725_ sky130_fd_sc_hd__o21bai_4
X_18763_ _09478_ _09479_ _09487_ VGND VGND VPWR VPWR _09652_ sky130_fd_sc_hd__a21oi_1
X_15975_ _06812_ _06849_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__and2_1
X_11098_ _02041_ _02040_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__nor2_4
X_17714_ _08575_ _08576_ _08561_ VGND VGND VPWR VPWR _08577_ sky130_fd_sc_hd__a21oi_2
XFILLER_76_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18694_ _09572_ _09574_ _09414_ _09415_ VGND VGND VPWR VPWR _09577_ sky130_fd_sc_hd__o2bb2ai_1
X_14926_ net739 net733 net663 net655 VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__nand4_2
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17645_ _08501_ _08503_ _08488_ VGND VGND VPWR VPWR _08509_ sky130_fd_sc_hd__o21ai_2
X_14857_ net716 net1012 VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__nand2_1
X_17576_ _08437_ net596 _08436_ net472 VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_63_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14788_ _09264_ _09493_ _05683_ _05685_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__o211ai_1
X_13808_ _04708_ net689 net752 VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__nand3_1
X_16527_ net307 _07389_ _07399_ VGND VGND VPWR VPWR _07400_ sky130_fd_sc_hd__a21oi_1
X_13739_ net393 _04642_ _04627_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_34_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19315_ _00483_ _10064_ net850 _00485_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__nand4_4
XFILLER_91_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16458_ _07195_ _07321_ _07328_ _07329_ VGND VGND VPWR VPWR _07331_ sky130_fd_sc_hd__o211ai_2
X_19246_ _10140_ _10141_ _10144_ VGND VGND VPWR VPWR _10146_ sky130_fd_sc_hd__nand3_1
X_16389_ net966 net950 net513 net506 VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__nand4_2
X_15409_ _06208_ _06209_ _06258_ _06260_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__and4_1
X_19177_ _10068_ _10063_ _10062_ VGND VGND VPWR VPWR _10071_ sky130_fd_sc_hd__nand3_4
XFILLER_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18128_ _09155_ _09210_ _09242_ _08970_ _08969_ VGND VGND VPWR VPWR _08976_ sky130_fd_sc_hd__o221ai_4
XFILLER_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18059_ _08905_ _08906_ VGND VGND VPWR VPWR _08908_ sky130_fd_sc_hd__nand2_1
XFILLER_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20021_ _01121_ _01137_ _01241_ _01243_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__o22ai_1
XFILLER_100_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer10 net806 VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer21 b_l\[1\] VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer43 a_l\[2\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 b_h\[10\] VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer54 _10059_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer76 net654 VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer87 b_h\[11\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer65 net861 VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer98 net894 VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_23_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20785_ clknet_leaf_26_clk _00425_ VGND VGND VPWR VPWR a_l\[7\] sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_12_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer100 net610 VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__buf_6
Xrebuffer111 net907 VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer133 net929 VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer155 _02669_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__buf_1
Xrebuffer144 a_l\[8\] VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__buf_2
XFILLER_108_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer177 a_l\[0\] VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer188 _03283_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__buf_1
Xrebuffer199 a_h\[12\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold570 term_high\[51\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12070_ _03002_ _03003_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__nand2_1
XFILLER_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11021_ _01961_ _01963_ _01958_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__nand3_1
XFILLER_89_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20219_ net727 net724 net551 net548 VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__nand4_1
XFILLER_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15760_ _06634_ _06636_ _06508_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__a21o_1
X_12972_ net659 net478 _03892_ _03895_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__a22o_1
X_11923_ _02753_ _02719_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__nand2_1
X_15691_ _06459_ _06499_ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__or2_1
XFILLER_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14711_ net730 net677 VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__nand2_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11854_ _02586_ _02592_ _02585_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__a21boi_2
XFILLER_122_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17430_ _08222_ _08292_ _08294_ VGND VGND VPWR VPWR _08296_ sky130_fd_sc_hd__nand3_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14642_ _05468_ _05471_ _05495_ _05542_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_103_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ net795 _01825_ _01826_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_45_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11785_ net653 net526 VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__nand2_1
X_17361_ _08222_ _08223_ net550 net516 VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__nand4_2
X_19100_ _09868_ _09988_ _09990_ VGND VGND VPWR VPWR _09991_ sky130_fd_sc_hd__nand3_4
X_14573_ _05471_ _05473_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__nor2_1
X_16312_ _07060_ _07182_ _07180_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__a21o_1
X_17292_ _08151_ _08157_ _08156_ VGND VGND VPWR VPWR _08160_ sky130_fd_sc_hd__o21ai_1
X_10736_ p_hl\[18\] p_lh\[18\] VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__and2_1
X_13524_ _04431_ _04399_ _04430_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__nand3_4
XFILLER_40_171 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16243_ net587 net561 net1063 net521 _07110_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__a41o_1
X_10667_ net794 _01707_ _01708_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__and3_1
X_13455_ _04335_ _04362_ _04363_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__nand3_4
X_19031_ _09919_ _09920_ VGND VGND VPWR VPWR _09922_ sky130_fd_sc_hd__nand2_1
X_16174_ _06950_ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__nand2_1
XFILLER_127_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ _03331_ _03332_ _03333_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__nand3_2
XFILLER_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10598_ _09690_ net1168 VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__and2_1
X_13386_ _04275_ _04277_ _04294_ _04295_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__o211ai_2
X_15125_ net733 net651 net911 net739 VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__a22oi_2
Xoutput108 net108 VGND VGND VPWR VPWR p[48] sky130_fd_sc_hd__buf_2
Xoutput119 net119 VGND VGND VPWR VPWR p[58] sky130_fd_sc_hd__buf_2
X_12337_ _03256_ _03266_ _03267_ _03269_ _03253_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__a32oi_2
XFILLER_56_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12268_ _02985_ _03173_ _03199_ _03200_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__o211ai_4
X_19933_ _00997_ _01041_ _01043_ _00998_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__a31o_1
X_15056_ _05938_ _05949_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__nand2_1
X_11219_ _02160_ _02158_ _02154_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_56_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19864_ _01079_ _01080_ VGND VGND VPWR VPWR _01081_ sky130_fd_sc_hd__nand2_1
X_14007_ _04912_ _04873_ _04911_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__nand3_4
X_12199_ net665 net501 VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__nand2_1
X_18815_ _09702_ _09704_ net231 VGND VGND VPWR VPWR _09708_ sky130_fd_sc_hd__nand3_4
Xoutput90 net90 VGND VGND VPWR VPWR p[31] sky130_fd_sc_hd__buf_2
X_19795_ net589 net580 net729 net725 VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_39_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15958_ _06832_ _06835_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__nand2_4
XFILLER_76_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18746_ _09546_ _09549_ _09626_ _09627_ VGND VGND VPWR VPWR _09633_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_39_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18677_ _09552_ _09554_ _09412_ VGND VGND VPWR VPWR _09558_ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_19_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14909_ _05446_ _05674_ _05801_ _05803_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__o22ai_4
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15889_ _06765_ _06766_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__nand2_1
X_17628_ net555 net500 net494 net560 VGND VGND VPWR VPWR _08492_ sky130_fd_sc_hd__a22oi_1
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17559_ _08414_ _08420_ _08419_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__o21a_1
X_20570_ clknet_leaf_29_clk _00210_ VGND VGND VPWR VPWR p_hh_pipe\[0\] sky130_fd_sc_hd__dfxtp_1
X_19229_ net1128 net717 _10124_ net216 VGND VGND VPWR VPWR _10128_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_118_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20004_ _01226_ _01227_ _01231_ VGND VGND VPWR VPWR _01232_ sky130_fd_sc_hd__nand3_2
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ _02498_ _02499_ _02496_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20768_ clknet_leaf_59_clk _00408_ VGND VGND VPWR VPWR a_h\[6\] sky130_fd_sc_hd__dfxtp_4
X_10521_ _01665_ _01668_ _01667_ net793 VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__o211a_1
XFILLER_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20699_ clknet_leaf_38_clk _00339_ VGND VGND VPWR VPWR p_lh\[1\] sky130_fd_sc_hd__dfxtp_1
X_13240_ _04143_ _04154_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__nand2_1
X_10452_ _01595_ _01616_ _01615_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__a21o_1
X_10383_ term_mid\[33\] term_high\[33\] _01557_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_131_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13171_ net890 _04092_ net138 VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_131_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12122_ _03053_ _03055_ _03050_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__a21o_1
X_16930_ net376 _07795_ _07798_ _07790_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__o211a_1
X_12053_ _02973_ _02981_ _02982_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__nand3_1
X_11004_ _01909_ _01946_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__nand2_1
XFILLER_104_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16861_ _07584_ _07586_ _07731_ net796 VGND VGND VPWR VPWR _07732_ sky130_fd_sc_hd__a31o_1
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15812_ _06676_ _06685_ _06686_ VGND VGND VPWR VPWR _06691_ sky130_fd_sc_hd__nand3_2
X_16792_ _07659_ _07661_ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__nor2_1
X_18600_ _09365_ _09380_ _09381_ _09237_ VGND VGND VPWR VPWR _09474_ sky130_fd_sc_hd__o2bb2ai_4
X_19580_ net1074 _00775_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__nand2_1
X_15743_ _06622_ _06585_ _06621_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__and3_4
X_18531_ _09394_ _09350_ VGND VGND VPWR VPWR _09399_ sky130_fd_sc_hd__nand2_1
X_12955_ _03880_ _03850_ _03844_ VGND VGND VPWR VPWR _03882_ sky130_fd_sc_hd__nand3b_2
XFILLER_46_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_5_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _09417_ _09646_ _02772_ _02836_ _02835_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__o221ai_4
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15674_ _06514_ _06547_ _06548_ VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__nand3_1
X_18462_ net252 _09296_ _09295_ _09290_ VGND VGND VPWR VPWR _09323_ sky130_fd_sc_hd__o2bb2ai_1
X_12886_ _03812_ _03813_ net669 net478 VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__and4_1
XFILLER_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11837_ net687 net492 VGND VGND VPWR VPWR _02774_ sky130_fd_sc_hd__nand2_1
X_17413_ _08277_ _08279_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__nand2_1
X_18393_ net604 net764 VGND VGND VPWR VPWR _09248_ sky130_fd_sc_hd__nand2_1
X_14625_ _05523_ _05524_ _05526_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__a21oi_1
X_11768_ net672 net511 VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__nand2_1
X_17344_ _08055_ _08207_ _08210_ _08052_ VGND VGND VPWR VPWR _08211_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_44_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _05289_ _05438_ _05454_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__nand3_4
XFILLER_147_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10719_ _01744_ _01748_ _01747_ p_hl\[14\] p_lh\[14\] VGND VGND VPWR VPWR _01752_
+ sky130_fd_sc_hd__a32o_1
X_13507_ net1058 net785 net673 net666 VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__nand4_2
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11699_ net462 _02636_ _02635_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__o21ai_1
X_17275_ _08138_ _08139_ _08040_ VGND VGND VPWR VPWR _08143_ sky130_fd_sc_hd__a21o_1
X_19014_ _09900_ _09901_ _09902_ _09759_ VGND VGND VPWR VPWR _09905_ sky130_fd_sc_hd__o2bb2ai_2
X_14487_ _05383_ _05385_ _05379_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__a21oi_1
Xrebuffer1 a_l\[3\] VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__clkbuf_2
X_16226_ net583 net572 net528 VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__nand3_1
X_13438_ net789 net673 VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nand2_2
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16157_ _07031_ net380 VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__or2_1
X_13369_ _04220_ _04223_ _04224_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_58_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16088_ _06898_ _06961_ net1127 net502 _06960_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__o2111ai_4
XFILLER_5_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15108_ _05950_ _05936_ _05937_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19916_ _01136_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__inv_2
X_15039_ _05931_ _05932_ _05924_ VGND VGND VPWR VPWR _05937_ sky130_fd_sc_hd__nand3_2
XFILLER_96_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19847_ _01061_ _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__and2_1
XFILLER_56_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19778_ _00744_ _00872_ _00871_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__o21ai_1
X_18729_ _09606_ _09608_ _09609_ VGND VGND VPWR VPWR _09615_ sky130_fd_sc_hd__a21o_1
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20622_ clknet_leaf_43_clk _00262_ VGND VGND VPWR VPWR p_ll_pipe\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20553_ clknet_leaf_26_clk _00193_ VGND VGND VPWR VPWR mid_sum\[16\] sky130_fd_sc_hd__dfxtp_1
X_20484_ clknet_leaf_45_clk _00124_ VGND VGND VPWR VPWR term_mid\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_105_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _03660_ _03662_ _03663_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__nand3_1
X_12671_ _03600_ _03601_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__nand2_1
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11622_ _02555_ _02557_ _02446_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15390_ net716 net657 _06281_ _06282_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__a22oi_4
X_14410_ _05308_ _05310_ _05299_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand3_2
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _05244_ _05118_ _05243_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__nand3_4
X_11553_ _02487_ _02488_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__nand2_2
X_10504_ net1320 _01656_ _01658_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__o21a_1
X_11484_ _02417_ _02421_ _02418_ VGND VGND VPWR VPWR _02424_ sky130_fd_sc_hd__nand3_4
X_17060_ _07781_ _07925_ net578 net503 _07924_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__o2111ai_1
X_14272_ _05172_ _05173_ _05145_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__a21oi_1
X_10435_ _01597_ _01598_ _01600_ _01602_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__o31a_1
X_16011_ _06874_ _06875_ net381 _06886_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__o2bb2ai_4
X_13223_ _04138_ net713 net777 _04137_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__and4_1
XFILLER_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13154_ net641 net634 net999 b_h\[14\] VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__nand4_1
X_12105_ a_h\[3\] net481 VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__nand2_1
XFILLER_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10366_ _01386_ _01375_ net797 VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a21oi_1
XFILLER_105_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17962_ net779 net632 _08813_ _08814_ VGND VGND VPWR VPWR _08815_ sky130_fd_sc_hd__a211o_1
X_13085_ _03969_ _03968_ _03963_ net394 VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__a22o_1
X_10297_ _00611_ _00622_ _00536_ _00569_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__o211ai_1
X_12036_ _02917_ _02969_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__nand2_1
X_17893_ _08723_ _08750_ _08722_ VGND VGND VPWR VPWR _08752_ sky130_fd_sc_hd__and3_1
X_16913_ _07671_ _07781_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_53_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19701_ net598 net718 VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__nand2_1
X_16844_ _07710_ _07711_ _07705_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__o21ai_1
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19632_ _00818_ _00825_ _00823_ _00780_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__o211ai_1
XFILLER_38_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16775_ net558 net554 b_h\[2\] net530 VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__and4_1
X_19563_ _00750_ _00751_ _00739_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__a21oi_1
X_13987_ net788 net643 VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__nand2_1
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15726_ net1090 net607 net531 net527 VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__and4_1
X_12938_ _03865_ _03796_ _03864_ VGND VGND VPWR VPWR _03866_ sky130_fd_sc_hd__nand3_1
X_18514_ _09237_ _09366_ _09376_ _09377_ VGND VGND VPWR VPWR _09380_ sky130_fd_sc_hd__o211ai_4
XFILLER_46_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _00681_ _00682_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__nand2_1
X_15657_ _09231_ _09526_ _06536_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__o21a_4
X_18445_ _09302_ _09215_ _09301_ VGND VGND VPWR VPWR _09305_ sky130_fd_sc_hd__and3_1
XFILLER_61_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12869_ _03736_ _03739_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__nor2_1
X_14608_ _05334_ net390 _05361_ _05368_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__o2bb2ai_2
X_15588_ _06466_ _06469_ _06463_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__a21o_1
X_18376_ _09161_ _09164_ VGND VGND VPWR VPWR _09229_ sky130_fd_sc_hd__nand2_1
X_17327_ _08176_ _08188_ _08191_ _08187_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__o211a_1
X_14539_ net761 net649 VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__nand2_1
X_17258_ _08124_ _08090_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__nand2_1
X_16209_ _06967_ _07063_ _07082_ _07083_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__o211ai_4
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17189_ net561 net559 net964 net969 VGND VGND VPWR VPWR _08057_ sky130_fd_sc_hd__nand4_4
XFILLER_143_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20605_ clknet_leaf_33_clk _00245_ VGND VGND VPWR VPWR p_ll_pipe\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20536_ clknet_leaf_45_clk _00176_ VGND VGND VPWR VPWR term_low\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20467_ clknet_leaf_14_clk _00107_ VGND VGND VPWR VPWR term_high\[59\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ net905 VGND VGND VPWR VPWR _09581_ sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_95_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20398_ clknet_leaf_46_clk _00038_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13910_ _04811_ _04813_ _04670_ net286 VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14890_ _05784_ _05786_ _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_126_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13841_ _02502_ _04134_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__nor2_2
X_16560_ _07428_ _07429_ _07431_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__o21bai_4
X_10984_ _01927_ _01928_ _01914_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__a21bo_1
XFILLER_74_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13772_ _04487_ _04550_ _04584_ _04678_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__o2111a_1
X_12723_ _03644_ _03649_ _03645_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__nand3_2
X_15511_ _06397_ _06399_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__nor2_1
X_16491_ _07361_ _07360_ _07359_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__nand3_2
X_18230_ _09075_ _09057_ VGND VGND VPWR VPWR _09077_ sky130_fd_sc_hd__nand2_1
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12654_ _03582_ _03583_ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a21bo_1
X_15442_ _06309_ _06331_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__xnor2_1
XFILLER_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11605_ _02519_ _02521_ _02536_ _02538_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18161_ _09002_ _08961_ VGND VGND VPWR VPWR _09009_ sky130_fd_sc_hd__nand2_1
X_12585_ _03261_ _03430_ _03433_ _03429_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__a22oi_4
X_15373_ net726 net640 VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__nand2_1
XFILLER_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11536_ _02473_ _02474_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__nand2_2
X_17112_ _07634_ _07789_ _07803_ _07979_ VGND VGND VPWR VPWR _07981_ sky130_fd_sc_hd__o211ai_2
X_18092_ _08938_ _08935_ _08899_ VGND VGND VPWR VPWR _08941_ sky130_fd_sc_hd__and3_1
X_14324_ _05223_ _05224_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__and3_1
XFILLER_144_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17043_ _07817_ _07909_ _07910_ VGND VGND VPWR VPWR _07912_ sky130_fd_sc_hd__nand3_2
Xwire352 _04450_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14255_ net788 net636 VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__nand2_1
X_11467_ _02401_ _02392_ _02400_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__nand3_2
XFILLER_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ _04094_ _04125_ _04123_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o21ai_1
X_10418_ net793 _01586_ _01587_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__and3_1
X_11398_ net1022 net495 VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__nand2_8
X_14186_ _05090_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__inv_2
XFILLER_112_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13137_ _04022_ _04019_ _04058_ _04057_ VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__a22oi_1
X_10349_ _01192_ _01203_ VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__nor2_1
X_18994_ _09882_ _09883_ VGND VGND VPWR VPWR _09885_ sky130_fd_sc_hd__nand2_4
XFILLER_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17945_ _08769_ _08788_ _08789_ VGND VGND VPWR VPWR _08802_ sky130_fd_sc_hd__o21a_1
X_13068_ _03990_ _03991_ _03992_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a21o_1
X_12019_ _02822_ _02947_ _02948_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__nand3_2
X_17876_ _08694_ _08698_ _08732_ _08734_ VGND VGND VPWR VPWR _08736_ sky130_fd_sc_hd__a22oi_1
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16827_ _07696_ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__nand2_1
Xclone264 net679 VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__clkbuf_16
XFILLER_65_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19615_ _00790_ _00792_ _00812_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__o21ai_2
XFILLER_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16758_ _07544_ _07542_ _07509_ _07547_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__a22oi_4
XFILLER_81_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19546_ _10170_ _00637_ _00639_ _00636_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__a22oi_4
X_15709_ net595 net542 VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_66_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16689_ _07486_ _07488_ _07555_ _07557_ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__nand4_1
XFILLER_22_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19477_ _00460_ _00461_ _00457_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18428_ _09282_ _09283_ _09267_ VGND VGND VPWR VPWR _09287_ sky130_fd_sc_hd__and3_1
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18359_ _09103_ _09109_ _09209_ net794 VGND VGND VPWR VPWR _09212_ sky130_fd_sc_hd__o31a_1
XFILLER_147_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20321_ net793 net18 VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__and2_1
XFILLER_128_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap652 net653 VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__buf_12
X_20252_ _01345_ _01404_ _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__nor3_1
Xmax_cap663 a_h\[10\] VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__buf_6
Xmax_cap641 a_h\[14\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_110_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap674 a_h\[8\] VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__buf_12
Xmax_cap696 a_h\[4\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__buf_8
Xmax_cap685 a_h\[6\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkbuf_8
X_20183_ net329 _01419_ _01422_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__a21oi_1
XFILLER_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12370_ _03175_ _03300_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_97_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11321_ _09395_ _09613_ _02190_ _02255_ _02258_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_97_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20519_ clknet_leaf_42_clk _00159_ VGND VGND VPWR VPWR term_low\[14\] sky130_fd_sc_hd__dfxtp_1
X_11252_ net706 net698 net510 net507 VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__nand4_2
X_14040_ _04917_ _04938_ _04768_ _04870_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_134_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11183_ _02120_ _02121_ _02125_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__nand3_4
XFILLER_121_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10203_ a_h\[2\] VGND VGND VPWR VPWR _09395_ sky130_fd_sc_hd__inv_6
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15991_ _06440_ _06867_ VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17730_ _08591_ _08592_ VGND VGND VPWR VPWR _08593_ sky130_fd_sc_hd__nand2_1
XFILLER_48_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14942_ _09362_ _09439_ _05836_ _05838_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_141_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ _08520_ _08522_ _08425_ VGND VGND VPWR VPWR _08525_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14873_ _05543_ _05547_ _05769_ _05770_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__o211ai_2
X_16612_ _07454_ _07479_ _07480_ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__nand3_1
X_13824_ net771 net667 VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__nand2_1
X_19400_ _00524_ _00526_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_106_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17592_ _08452_ _08455_ _08372_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__nand3_2
X_19331_ net887 net603 _05043_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__and3_1
X_16543_ _07350_ _07412_ _07413_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__nand3_4
X_10967_ _01910_ net466 _01907_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o21bai_4
XTAP_TAPCELL_ROW_106_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ net734 net1077 net703 net741 VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__a22o_1
XFILLER_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16474_ _07344_ _07346_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__nand2_1
X_12706_ net659 net490 VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__nand2_1
X_13686_ net789 net656 VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__nand2_1
X_10898_ net794 net1330 VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__and2_1
X_19262_ net1086 net552 _09155_ VGND VGND VPWR VPWR _10163_ sky130_fd_sc_hd__a21o_1
X_18213_ _09242_ _08970_ _08965_ _08968_ VGND VGND VPWR VPWR _09060_ sky130_fd_sc_hd__o22ai_2
X_12637_ _03563_ _03565_ _03566_ VGND VGND VPWR VPWR _03568_ sky130_fd_sc_hd__a21o_1
X_19193_ net598 net592 net744 net738 VGND VGND VPWR VPWR _10089_ sky130_fd_sc_hd__nand4_4
X_15425_ _09351_ _09515_ _06266_ _06269_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_139_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18144_ _08983_ _08986_ _08988_ VGND VGND VPWR VPWR _08992_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_61_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12568_ _03485_ net176 _03377_ _03483_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__o22a_1
X_15356_ _06247_ _06248_ _06240_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__and3_1
XFILLER_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11519_ _02455_ _02456_ _02452_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__a21o_1
X_18075_ net779 net611 _08920_ _08921_ VGND VGND VPWR VPWR _08924_ sky130_fd_sc_hd__a22o_1
X_12499_ net644 net511 net508 net1016 VGND VGND VPWR VPWR _03431_ sky130_fd_sc_hd__a22o_1
X_15287_ _06180_ _06172_ _06000_ _06181_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__o211ai_4
X_14307_ _09308_ _09417_ _05053_ _05207_ _05206_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__o221ai_2
Xwire193 _05269_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_2
X_17026_ _07893_ _07894_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__nand2_1
X_14238_ _05132_ _05135_ _05134_ _05120_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__o211ai_2
XFILLER_131_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14169_ _05068_ _05069_ _05040_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__nand3_1
XFILLER_140_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18977_ _09739_ _09852_ _09853_ VGND VGND VPWR VPWR _09868_ sky130_fd_sc_hd__a21boi_4
XFILLER_140_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17928_ _08784_ _08785_ VGND VGND VPWR VPWR _08786_ sky130_fd_sc_hd__nor2_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_0_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17859_ net937 net484 net480 net875 VGND VGND VPWR VPWR _08719_ sky130_fd_sc_hd__a22o_1
XFILLER_38_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_497 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_19529_ _00685_ _00694_ _00697_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__o21ai_1
XFILLER_62_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer304 _09918_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__buf_1
XFILLER_108_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer337 _04452_ VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__buf_2
Xrebuffer315 b_h\[13\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer326 net776 VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__buf_6
Xrebuffer348 _05163_ VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_146_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20304_ _01540_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__nor2_1
XFILLER_116_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap460 _03312_ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_92_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20235_ _01478_ _01475_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__nand2_1
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap471 _01268_ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_1
Xmax_cap493 net494 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20166_ _01345_ _01352_ _01404_ _01344_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__o211ai_1
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20097_ _01323_ _01329_ _01330_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__nand3_1
XFILLER_39_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11870_ _02698_ _02804_ _02803_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__and3_1
X_10821_ _01837_ _01832_ _01831_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__a21o_1
XFILLER_53_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10752_ p_hl\[19\] p_lh\[19\] p_hl\[18\] p_lh\[18\] VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__o211a_1
X_13540_ _04446_ _04447_ _04448_ _04341_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_71_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13471_ _04375_ _04376_ _04379_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__nand3_2
XFILLER_41_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12422_ _03346_ _03347_ _03352_ _03353_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10683_ _01716_ _01719_ _01720_ net797 VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__a31o_1
XFILLER_13_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15210_ _06101_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__nor2_2
X_16190_ _02338_ _06441_ _07026_ _07027_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__o22ai_2
XFILLER_138_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12353_ _02899_ _02996_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__o21ai_4
X_15141_ _06026_ _06030_ _06033_ _06015_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_134_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11304_ net361 _02205_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__and2_1
X_12284_ _03125_ _03214_ _03215_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__nand3_2
XFILLER_107_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15072_ _05819_ _05903_ _05965_ _05966_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__a22o_1
X_11235_ _02088_ _02080_ _02172_ _02173_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__o211ai_4
X_18900_ _09786_ _09787_ _09788_ VGND VGND VPWR VPWR _09792_ sky130_fd_sc_hd__nand3_1
X_14023_ _09264_ _09428_ _04927_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__o21ai_2
XFILLER_122_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19880_ _00872_ _00982_ _00987_ VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__o21a_1
X_11166_ net712 net501 VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__nand2_1
X_18831_ net275 _09572_ _09573_ net185 VGND VGND VPWR VPWR _09724_ sky130_fd_sc_hd__o2bb2ai_2
X_15974_ net260 VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__inv_2
X_11097_ _01944_ _01948_ _01947_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__o21a_1
XFILLER_110_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18762_ _09642_ _09649_ _09650_ VGND VGND VPWR VPWR _09651_ sky130_fd_sc_hd__o21ai_2
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17713_ _08569_ _08572_ _08573_ VGND VGND VPWR VPWR _08576_ sky130_fd_sc_hd__nand3_4
XFILLER_0_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14925_ _05821_ _05822_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__nand2_1
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18693_ net185 _09573_ _09572_ net275 VGND VGND VPWR VPWR _09576_ sky130_fd_sc_hd__o211ai_2
X_17644_ _08488_ _08502_ _08504_ VGND VGND VPWR VPWR _08508_ sky130_fd_sc_hd__nand3b_1
X_14856_ _05755_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__inv_2
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17575_ _08436_ _08437_ _08432_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_63_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14787_ _05683_ _05685_ net745 net655 VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__nand4_2
X_13807_ _04632_ _04707_ net746 net694 _04711_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__o2111ai_4
X_11999_ _02858_ _02929_ _02824_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__a21o_1
X_16526_ _07391_ _07395_ _07398_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__o21ai_4
X_13738_ _04628_ net393 _04642_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_34_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19314_ _10058_ _10064_ _00483_ _00485_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__and4_1
X_19245_ _10140_ _10141_ _10144_ VGND VGND VPWR VPWR _10145_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_14_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16457_ _07195_ _07321_ _07328_ _07329_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__o211a_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13669_ _04466_ _04473_ _04576_ _04577_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o211ai_2
X_16388_ a_l\[7\] net506 VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__nand2_1
X_15408_ _06299_ _06300_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__nand2_1
X_19176_ _10066_ _10067_ _10065_ VGND VGND VPWR VPWR _10070_ sky130_fd_sc_hd__nand3_4
X_18127_ _08969_ _08971_ _08965_ VGND VGND VPWR VPWR _08975_ sky130_fd_sc_hd__a21o_1
X_15339_ _06165_ _06161_ _06163_ _06232_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__o211ai_4
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18058_ net615 net774 net769 net623 VGND VGND VPWR VPWR _08907_ sky130_fd_sc_hd__a22oi_1
XFILLER_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17009_ _07878_ _07872_ _07873_ VGND VGND VPWR VPWR _07879_ sky130_fd_sc_hd__nand3_2
XFILLER_99_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20020_ net332 _01136_ _01242_ _01244_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__nand4_1
XFILLER_140_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer11 b_l\[4\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer44 a_l\[2\] VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer33 b_h\[10\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer55 _09889_ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer22 b_l\[7\] VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer77 a_l\[14\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__buf_2
Xrebuffer88 net884 VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__buf_2
Xrebuffer66 net861 VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer99 b_l\[8\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd1_1
X_20784_ clknet_leaf_26_clk _00424_ VGND VGND VPWR VPWR a_l\[6\] sky130_fd_sc_hd__dfxtp_4
Xrebuffer112 net907 VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer101 _10019_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__buf_6
Xrebuffer156 net766 VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__buf_6
Xrebuffer123 net669 VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__buf_2
Xrebuffer145 net941 VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer134 _05177_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__buf_6
Xrebuffer189 net688 VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__buf_2
Xhold560 _00072_ VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold571 term_low\[30\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ net691 net1106 _01961_ _01963_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__a22o_1
XFILLER_103_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap290 _03564_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__buf_1
XFILLER_2_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20218_ _01410_ _01459_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__nand2_1
X_20149_ _01284_ _01287_ _01315_ _01383_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__o211ai_2
XFILLER_58_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12971_ _03892_ _03895_ _03890_ VGND VGND VPWR VPWR _03898_ sky130_fd_sc_hd__a21oi_2
X_11922_ _02855_ _02857_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__nand2_2
X_15690_ _06568_ _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__nand2_1
X_14710_ _05478_ _05481_ _05480_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__a21boi_1
X_11853_ _02788_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__nand2_1
X_14641_ _05488_ _05492_ _05489_ _05496_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_103_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _01824_ _01821_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__nand2_1
X_17360_ _08223_ _08041_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_45_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _07059_ _07183_ _07185_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__a21oi_4
X_11784_ _02624_ _02638_ _02622_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__a21o_1
X_14572_ net720 net699 _05469_ _05470_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__a22o_1
X_17291_ _08151_ _08157_ _08156_ VGND VGND VPWR VPWR _08159_ sky130_fd_sc_hd__o21a_1
X_10735_ p_hl\[18\] p_lh\[18\] VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__nor2_1
X_13523_ _04409_ _04427_ _04428_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__nand3b_1
XFILLER_15_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16242_ _07114_ net515 net950 VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__and3_1
X_10666_ _01703_ _01704_ _01706_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__or3_1
X_13454_ _04361_ _04334_ _04360_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__nand3_1
X_19030_ _09917_ _09920_ VGND VGND VPWR VPWR _09921_ sky130_fd_sc_hd__nand2_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16173_ _07044_ _07046_ _06812_ _06849_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__o2bb2ai_1
X_12405_ _03331_ _03333_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__nand2_1
X_13385_ _04278_ _04279_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__o21ai_1
X_10597_ _09690_ net1163 VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__and2_1
X_15124_ net739 net733 net651 net911 VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__nand4_2
Xoutput109 net109 VGND VGND VPWR VPWR p[49] sky130_fd_sc_hd__buf_2
XFILLER_126_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12336_ _03264_ _03265_ _03255_ VGND VGND VPWR VPWR _03269_ sky130_fd_sc_hd__nand3_4
XPHY_EDGE_ROW_81_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12267_ _03193_ _03197_ _03174_ _03198_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__o211ai_4
X_19932_ _01153_ _01154_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__nand2_1
X_15055_ _05945_ _05947_ _05937_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__o21ai_1
X_11218_ net1078 net681 net525 net519 VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__nand4_2
X_12198_ net661 net653 net511 net508 VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_56_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19863_ _01077_ _01076_ _01075_ VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__nand3_2
X_14006_ _04884_ _04885_ _04903_ _04905_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__o22ai_2
Xoutput91 net91 VGND VGND VPWR VPWR p[32] sky130_fd_sc_hd__buf_2
XFILLER_122_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11149_ _02085_ net465 _02077_ _02084_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__o211ai_4
XFILLER_68_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18814_ _09511_ _09520_ _09705_ net217 VGND VGND VPWR VPWR _09707_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_56_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput80 net80 VGND VGND VPWR VPWR p[22] sky130_fd_sc_hd__buf_2
XFILLER_95_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19794_ net580 net729 VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15957_ _06829_ _06830_ _06741_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__nand3_2
XFILLER_83_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18745_ _09546_ _09549_ _09627_ _09626_ VGND VGND VPWR VPWR _09632_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15888_ _06760_ _06762_ _06756_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__a21o_1
XFILLER_64_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18676_ _09553_ _09555_ _09412_ VGND VGND VPWR VPWR _09557_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_19_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14908_ _05802_ _05804_ _05675_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_90_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17627_ net555 net500 VGND VGND VPWR VPWR _08491_ sky130_fd_sc_hd__nand2_1
XFILLER_63_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14839_ _05728_ _05734_ _05733_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__o21ai_2
X_17558_ _08413_ _08415_ _08418_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__a21o_1
X_16509_ _07231_ _07377_ net1004 net541 _07376_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__o2111ai_1
X_17489_ _08336_ _08340_ _08351_ _08350_ VGND VGND VPWR VPWR _08355_ sky130_fd_sc_hd__o211ai_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19228_ _09900_ _10123_ _10122_ VGND VGND VPWR VPWR _10127_ sky130_fd_sc_hd__a21oi_1
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19159_ _09220_ _09297_ _10044_ _10045_ VGND VGND VPWR VPWR _10052_ sky130_fd_sc_hd__o211ai_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_141_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20003_ _01114_ _01122_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nand2_1
XFILLER_140_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_129_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20767_ clknet_leaf_59_clk _00407_ VGND VGND VPWR VPWR a_h\[5\] sky130_fd_sc_hd__dfxtp_4
X_10520_ _01665_ _01668_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__nor2_2
X_10451_ net443 _01599_ _01603_ _01609_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_138_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20698_ clknet_leaf_38_clk _00338_ VGND VGND VPWR VPWR p_lh\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10382_ term_mid\[32\] term_high\[32\] term_mid\[33\] term_high\[33\] VGND VGND VPWR
+ VPWR _01557_ sky130_fd_sc_hd__a22o_1
X_13170_ net853 _04092_ net138 VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_131_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12121_ _02836_ _03051_ _03050_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__o21ai_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold390 mid_sum\[21\] VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12052_ _02983_ _02984_ _02972_ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__a21oi_1
XFILLER_78_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11003_ net697 net1109 net1052 net702 VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__a22oi_1
XFILLER_78_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16860_ _07726_ _07729_ _07728_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o21a_1
X_15811_ _06599_ _06606_ _06686_ _06604_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__o211ai_1
X_16791_ _07633_ _07635_ _07657_ VGND VGND VPWR VPWR _07662_ sky130_fd_sc_hd__o21ai_1
X_15742_ _06617_ _06596_ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__nand2_1
X_18530_ net303 _09347_ _09394_ VGND VGND VPWR VPWR _09398_ sky130_fd_sc_hd__o21ai_2
X_12954_ _03843_ _03849_ _03880_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__o21ai_4
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _02835_ _02837_ _02838_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21o_1
X_18461_ net153 _09312_ _09315_ _09320_ VGND VGND VPWR VPWR _09322_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15673_ _06550_ _06551_ _06513_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__a21oi_4
X_17412_ _08156_ _08272_ _08274_ _08027_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__a22oi_1
XFILLER_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12885_ net659 net654 b_h\[12\] b_h\[13\] VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__nand4_1
X_11836_ _02771_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__nand2_1
X_18392_ _09244_ _09245_ _09232_ VGND VGND VPWR VPWR _09247_ sky130_fd_sc_hd__nand3_2
XFILLER_61_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14624_ b_l\[15\] net709 _05385_ _05384_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__a31o_1
X_11767_ net682 net501 VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__nand2_1
X_17343_ net554 net969 VGND VGND VPWR VPWR _08210_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_44_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14555_ net1000 _05291_ _05452_ _05453_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__a22oi_1
X_17274_ _08138_ _08139_ _08040_ VGND VGND VPWR VPWR _08142_ sky130_fd_sc_hd__a21oi_1
X_10718_ p_hl\[15\] p_lh\[15\] VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__xor2_1
X_13506_ net785 net666 VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_24_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11698_ _09460_ _09602_ _02630_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o21ai_1
X_16225_ net582 net573 VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__nand2_4
X_19013_ _09760_ _09900_ _09901_ _09903_ VGND VGND VPWR VPWR _09904_ sky130_fd_sc_hd__nand4_2
X_14486_ _05379_ _05383_ _05385_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__and3_1
Xrebuffer2 net798 VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd1_1
X_10649_ p_hl\[4\] p_lh\[4\] VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__nand2_1
X_13437_ net777 net932 VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__nand2_1
X_16156_ _06847_ _07029_ net422 VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__nor3_2
XFILLER_115_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13368_ _04274_ _04276_ _04275_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_58_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16087_ net1127 net502 _06960_ _06962_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__a22o_1
X_12319_ _03125_ _03214_ _03215_ _03219_ _03231_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__a32oi_2
XFILLER_114_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15107_ _06002_ net945 VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13299_ _04211_ _04212_ _09690_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__and3_1
X_19915_ _01132_ _01133_ _01124_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__o21ai_2
X_15038_ _05931_ _05932_ _05924_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__a21oi_2
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19846_ _01060_ net598 _01059_ net717 VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__nand4_2
X_16989_ net845 net472 _07856_ _07857_ VGND VGND VPWR VPWR _07859_ sky130_fd_sc_hd__a22o_1
X_19777_ _00983_ _00984_ _00981_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__nand3_2
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18728_ _09606_ _09608_ _09609_ VGND VGND VPWR VPWR _09614_ sky130_fd_sc_hd__a21oi_2
XFILLER_36_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18659_ net621 net618 net743 net737 VGND VGND VPWR VPWR _09539_ sky130_fd_sc_hd__nand4_4
XFILLER_52_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20621_ clknet_leaf_43_clk _00261_ VGND VGND VPWR VPWR p_ll_pipe\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20552_ clknet_leaf_54_clk _00192_ VGND VGND VPWR VPWR mid_sum\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20483_ clknet_leaf_43_clk _00123_ VGND VGND VPWR VPWR term_mid\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12670_ _03486_ _03489_ _03597_ _03599_ VGND VGND VPWR VPWR _03601_ sky130_fd_sc_hd__nand4b_1
X_11621_ _02446_ _02555_ _02557_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__nand3_2
XFILLER_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14340_ _05186_ _05190_ _05232_ _05234_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__o2bb2ai_1
X_11552_ _02483_ _02489_ _02490_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10503_ _01653_ _01657_ net796 VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__a21oi_1
X_11483_ _02419_ _02420_ _02422_ VGND VGND VPWR VPWR _02423_ sky130_fd_sc_hd__nand3_2
Xwire534 b_h\[2\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__buf_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14271_ _05171_ _05155_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__nand2_1
X_10434_ net796 _01601_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__nor2_1
X_16010_ _06883_ _06884_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__nor2_1
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire578 a_l\[10\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__buf_12
X_13222_ _04137_ _04138_ _09155_ _09177_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__o2bb2a_1
X_13153_ net634 net999 b_h\[14\] net641 VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__a22o_1
X_10365_ net471 _01322_ net1369 VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__o21ai_1
X_12104_ net358 _02875_ _02873_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__a21boi_2
XFILLER_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17961_ net623 net790 net781 net627 VGND VGND VPWR VPWR _08814_ sky130_fd_sc_hd__a22oi_2
X_13084_ _04007_ _04000_ _04006_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__nand3b_2
X_10296_ _00536_ _00569_ _00611_ _00622_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__a211o_1
X_12035_ _02876_ _02878_ _02917_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__o21ai_1
X_17892_ _08723_ _08722_ _08750_ VGND VGND VPWR VPWR _08751_ sky130_fd_sc_hd__a21oi_1
X_16912_ net571 net513 net506 net1093 VGND VGND VPWR VPWR _07782_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_53_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19700_ _00899_ _00900_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__nand2_1
X_16843_ _07705_ _07712_ VGND VGND VPWR VPWR _07714_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19631_ _00777_ _00823_ _00826_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_144_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19562_ net445 _00755_ _00740_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__o21ai_2
X_16774_ net554 net530 VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__nand2_1
X_18513_ _09375_ net581 net780 VGND VGND VPWR VPWR _09379_ sky130_fd_sc_hd__nand3_1
X_13986_ net778 net656 VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__nand2_1
X_15725_ net612 net608 VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__nand2_8
X_12937_ _03804_ _03805_ _03857_ net175 VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19493_ _00677_ net298 _00678_ _00679_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__nand4_4
XFILLER_33_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15656_ net602 net1041 VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__nand2_4
X_18444_ _09184_ _09213_ _09299_ _09300_ VGND VGND VPWR VPWR _09304_ sky130_fd_sc_hd__o211ai_2
X_12868_ _03775_ _03725_ _03774_ VGND VGND VPWR VPWR _03796_ sky130_fd_sc_hd__o21ai_1
XFILLER_61_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11819_ _02753_ _02719_ _02752_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__nand3_1
X_18375_ _09161_ _09145_ VGND VGND VPWR VPWR _09228_ sky130_fd_sc_hd__nand2_1
X_14607_ net716 net703 VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__nand2_1
XFILLER_21_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15587_ net628 net607 net542 net522 VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__nand4_1
X_17326_ _08187_ _08189_ _08191_ VGND VGND VPWR VPWR _08193_ sky130_fd_sc_hd__a21o_1
X_12799_ net1049 net634 b_h\[7\] b_h\[8\] VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__and4_2
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14538_ _09220_ _09504_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__nor2_1
X_17257_ _08122_ _08092_ _08121_ _08091_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__a31oi_2
X_14469_ _05362_ _05368_ _05366_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__a21oi_1
X_16208_ _07074_ _07076_ _07078_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__a21o_1
X_17188_ net561 net1004 net964 net969 VGND VGND VPWR VPWR _08056_ sky130_fd_sc_hd__and4_1
XFILLER_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16139_ _07011_ _07013_ _06977_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__a21oi_1
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19829_ _01036_ _01037_ _01039_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__nand3_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20604_ clknet_leaf_35_clk _00244_ VGND VGND VPWR VPWR p_ll_pipe\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20535_ clknet_leaf_45_clk _00175_ VGND VGND VPWR VPWR term_low\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20466_ clknet_leaf_14_clk _00106_ VGND VGND VPWR VPWR term_high\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20397_ clknet_leaf_47_clk _00037_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13840_ _04744_ _04745_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__nand2_2
X_10983_ _01908_ _01912_ _01913_ _01927_ _01928_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__o2111ai_4
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13771_ _04655_ _04660_ _04673_ _04674_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__o2bb2ai_2
X_16490_ _07359_ _07360_ _07361_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12722_ _03646_ _03647_ _03650_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__nand3_2
X_15510_ net795 _06396_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__nand2_1
XFILLER_16_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_90_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15441_ _06292_ _06296_ _06331_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__and3_1
XFILLER_31_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12653_ _09428_ _09679_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__nor2_1
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11604_ _02519_ _02521_ _02537_ _02539_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__nand4_2
X_18160_ _09006_ _09000_ VGND VGND VPWR VPWR _09008_ sky130_fd_sc_hd__nand2_2
X_12584_ _03511_ _03512_ _03151_ _03420_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15372_ net722 net643 VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__nand2_1
X_11535_ _02347_ _02468_ _02470_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__nand3_1
X_17111_ _07963_ _07964_ _07974_ VGND VGND VPWR VPWR _07980_ sky130_fd_sc_hd__a21oi_2
X_18091_ _08935_ _08938_ _08899_ VGND VGND VPWR VPWR _08940_ sky130_fd_sc_hd__a21o_1
Xwire320 _04073_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__buf_1
X_14323_ _05050_ _05065_ _05063_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__o21ai_1
Xwire331 _01307_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__buf_1
XFILLER_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire364 _01863_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__buf_1
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17042_ _07909_ _07910_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__nand2_1
Xwire375 _08102_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_1
X_14254_ net778 net643 VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__nand2_2
Xwire386 _06581_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
X_11466_ _02402_ _02405_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__nand2_1
X_13205_ _04093_ _04124_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__nand2_1
Xwire397 _03731_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10417_ _01579_ _01583_ _01585_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__or3_1
X_11397_ _02248_ _02316_ _02315_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__a21boi_1
XFILLER_99_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14185_ _04837_ _05087_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__xor2_2
XFILLER_140_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13136_ _03960_ _03963_ _03975_ _09679_ _09493_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a311o_1
X_18993_ net1113 net1082 net737 net603 VGND VGND VPWR VPWR _09884_ sky130_fd_sc_hd__a22oi_4
X_10348_ term_low\[29\] term_mid\[29\] VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__nor2_1
X_17944_ _08769_ _08788_ VGND VGND VPWR VPWR _08801_ sky130_fd_sc_hd__nor2_1
X_13067_ _03990_ _03991_ _03992_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__a21oi_1
X_10279_ net1360 _10158_ _00450_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__o21a_1
X_12018_ _02947_ _02948_ _02822_ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__a21o_1
Xclone221 net511 VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__clkbuf_16
X_17875_ _08732_ _08734_ VGND VGND VPWR VPWR _08735_ sky130_fd_sc_hd__nand2_1
XFILLER_39_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16826_ net236 _07694_ _07629_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__nand3_4
Xclone265 net544 net540 VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__nand2_4
XFILLER_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19614_ _00793_ _00811_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__nand2_2
X_16757_ _07626_ _07627_ VGND VGND VPWR VPWR _07628_ sky130_fd_sc_hd__nand2_1
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclone287 net565 VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__clkbuf_16
X_19545_ net919 net552 net407 _00736_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__a31o_1
X_13969_ net771 net660 VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__nand2_1
X_15708_ net617 net522 VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16688_ _07486_ _07488_ _07555_ _07557_ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__and4_1
X_19476_ _00460_ _00461_ _00457_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__a21o_1
X_15639_ net612 net531 VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18427_ _09282_ _09283_ _09267_ VGND VGND VPWR VPWR _09285_ sky130_fd_sc_hd__a21o_1
X_18358_ _09106_ _09102_ _09104_ VGND VGND VPWR VPWR _09211_ sky130_fd_sc_hd__o21ai_1
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17309_ _08174_ net449 _08167_ _08175_ VGND VGND VPWR VPWR _08176_ sky130_fd_sc_hd__o211a_1
X_18289_ net774 net1113 VGND VGND VPWR VPWR _09135_ sky130_fd_sc_hd__nand2_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20320_ net793 net17 VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__and2_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap620 a_l\[3\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__buf_12
XFILLER_115_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap631 net632 VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__buf_6
Xmax_cap653 net654 VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__buf_12
X_20251_ _01490_ _01449_ _01448_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__nand3_1
Xmax_cap642 net643 VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_8
Xmax_cap697 net698 VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__buf_6
Xmax_cap686 net687 VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_110_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap664 net665 VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__buf_12
Xmax_cap675 net676 VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__buf_8
X_20182_ _01366_ _01421_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__nand2_1
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11320_ _02257_ _02258_ _02254_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_97_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20518_ clknet_leaf_41_clk _00158_ VGND VGND VPWR VPWR term_low\[13\] sky130_fd_sc_hd__dfxtp_1
X_20449_ clknet_leaf_17_clk _00089_ VGND VGND VPWR VPWR term_high\[41\] sky130_fd_sc_hd__dfxtp_1
X_11251_ net698 net507 VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__nand2_1
XFILLER_109_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11182_ _02035_ net363 _02033_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__a21oi_4
XFILLER_107_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ net715 VGND VGND VPWR VPWR _09384_ sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_128_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15990_ net594 net586 VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__nand2_8
XFILLER_79_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14941_ _05837_ _05839_ net720 net685 VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_141_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17660_ _08522_ _08425_ _08520_ VGND VGND VPWR VPWR _08524_ sky130_fd_sc_hd__nand3_2
XFILLER_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14872_ _05543_ _05547_ _05769_ _05770_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__o211a_1
X_16611_ _07482_ _07453_ _07481_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__nand3_2
X_17591_ _08451_ _08454_ _08372_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__o21bai_4
XFILLER_75_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13823_ net1122 net670 VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__nand2_1
X_16542_ _07410_ net255 _07351_ _07411_ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__o211ai_2
X_19330_ _00502_ _00503_ _00495_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__nand3_1
X_10966_ _09177_ _09602_ _01911_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__o21ai_4
XTAP_TAPCELL_ROW_106_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13754_ net734 net709 net703 net741 VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__a22oi_1
X_16473_ _07338_ _07341_ _07339_ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__nand3_1
X_12705_ net659 net490 VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__and2_1
X_13685_ net783 net660 VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__nand2_1
XFILLER_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10897_ net794 net1198 VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__and2_1
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19261_ _10040_ _10161_ VGND VGND VPWR VPWR _10162_ sky130_fd_sc_hd__nand2_2
X_18212_ _08965_ _08971_ VGND VGND VPWR VPWR _09059_ sky130_fd_sc_hd__nand2_1
X_12636_ _03563_ _03565_ _03566_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__a21oi_1
X_19192_ net592 net744 VGND VGND VPWR VPWR _10088_ sky130_fd_sc_hd__nand2_1
X_15424_ net388 _06315_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_139_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _08988_ net764 net623 _08986_ VGND VGND VPWR VPWR _08991_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_61_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _06247_ _06248_ _06240_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__a21oi_1
X_12567_ _03495_ _03497_ _03498_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__o21a_1
XFILLER_79_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire150 _06259_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_1
X_14306_ _05206_ _05208_ _09308_ _09417_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11518_ _01871_ _02338_ _02452_ _02456_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__o211ai_1
X_18074_ net459 _06681_ net779 net611 _08920_ VGND VGND VPWR VPWR _08923_ sky130_fd_sc_hd__o2111ai_1
X_12498_ net644 net514 VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__nand2_2
X_15286_ _06173_ _06175_ _06158_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__a21o_1
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11449_ _02383_ _02384_ net327 VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__nand3_4
X_17025_ _07890_ _07892_ _07887_ VGND VGND VPWR VPWR _07894_ sky130_fd_sc_hd__nand3b_1
X_14237_ _05134_ _05136_ _05120_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__and3_1
XFILLER_131_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14168_ _05070_ _05064_ _05041_ _05071_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__o211ai_4
XFILLER_98_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13119_ net634 net1151 net999 net641 VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a22o_1
X_18976_ _09850_ net832 _09866_ VGND VGND VPWR VPWR _09867_ sky130_fd_sc_hd__o21ai_1
X_14099_ _04972_ _05002_ _05003_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__nand3_2
X_17927_ _09373_ _09668_ _08781_ _08783_ _08758_ VGND VGND VPWR VPWR _08785_ sky130_fd_sc_hd__o311a_1
X_17858_ net874 net936 net484 net480 VGND VGND VPWR VPWR _08718_ sky130_fd_sc_hd__nand4_1
XFILLER_78_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16809_ _07666_ _07673_ _07675_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__and3_1
XFILLER_94_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17789_ _08586_ _08650_ _08648_ VGND VGND VPWR VPWR _08651_ sky130_fd_sc_hd__and3_1
X_19528_ net183 _00718_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19459_ net1074 VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__inv_2
XFILLER_147_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer327 net1123 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_79_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20303_ _01521_ _01539_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__nor2_1
XFILLER_146_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap461 _03052_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_2
XFILLER_104_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap450 _08095_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_2
XFILLER_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap472 net473 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_6
X_20234_ _01469_ _01472_ _01473_ _01468_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__a31oi_1
XFILLER_115_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap494 net495 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__buf_12
X_20165_ _01344_ _01355_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_110_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20096_ _01329_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__nand2_1
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_84_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10820_ p_hl\[29\] net1361 VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__xor2_1
XFILLER_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10751_ _01777_ _01778_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__nor2_1
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13470_ _04377_ _04378_ _04380_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__nand3_1
XFILLER_139_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12421_ _03352_ _03353_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__nand2_1
X_10682_ _01716_ _01719_ _01720_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__a21oi_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ _03283_ _03284_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__nor2_2
X_15140_ _05913_ _06035_ _06036_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__nand3_2
X_11303_ _02242_ _02243_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__or2_1
XFILLER_126_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12283_ _03169_ _03171_ _03205_ _03207_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__o2bb2ai_1
X_15071_ _05819_ _05903_ _05965_ _05966_ VGND VGND VPWR VPWR _05969_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_134_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11234_ _02175_ _02164_ _02174_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__nand3_4
XFILLER_5_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14022_ _04708_ _04925_ net746 net689 _04924_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__o2111ai_4
XFILLER_136_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11165_ net707 net702 net510 net507 VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__nand4_2
XFILLER_122_654 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18830_ _09572_ net275 VGND VGND VPWR VPWR _09723_ sky130_fd_sc_hd__nand2_1
X_15973_ _06812_ _06849_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__nor2_1
X_11096_ _02038_ _02039_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__or2_4
XFILLER_121_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18761_ net763 net943 _09643_ _09645_ VGND VGND VPWR VPWR _09650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17712_ _08568_ _08571_ _08573_ VGND VGND VPWR VPWR _08575_ sky130_fd_sc_hd__o21bai_4
X_14924_ net733 net662 net655 net739 VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__a22oi_4
X_18692_ net185 _09573_ _09572_ VGND VGND VPWR VPWR _09575_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17643_ _08486_ _08487_ _08502_ _08504_ VGND VGND VPWR VPWR _08507_ sky130_fd_sc_hd__and4_1
XFILLER_48_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14855_ _05467_ _05604_ net389 _05629_ _05634_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__o2111ai_4
XFILLER_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11998_ _02929_ _02858_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__nand2_1
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17574_ net596 net472 _08436_ _08437_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__a22o_1
XFILLER_63_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14786_ _05683_ _05685_ _05680_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__a21bo_1
XFILLER_35_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13806_ _04710_ _04711_ _04706_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a21o_1
X_10949_ _01892_ _01893_ _01894_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__a21o_1
X_16525_ _07391_ _07393_ _07390_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__o21bai_2
XFILLER_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13737_ _04628_ net393 _04642_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__and3_1
XFILLER_32_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19313_ _00481_ _00480_ net851 _00487_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__nand4_4
X_16456_ _07324_ _07326_ _09188_ _09646_ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__o2bb2ai_2
X_19244_ _09166_ _09384_ _09980_ _09979_ VGND VGND VPWR VPWR _10144_ sky130_fd_sc_hd__o31a_2
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13668_ _04570_ _04572_ _04393_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__o21bai_4
X_15407_ _06297_ _06257_ _06254_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_14_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16387_ _07131_ _07260_ VGND VGND VPWR VPWR _07261_ sky130_fd_sc_hd__nand2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12619_ net674 net483 VGND VGND VPWR VPWR _03550_ sky130_fd_sc_hd__nand2_1
X_13599_ net924 net768 net683 net675 VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__nand4_4
X_19175_ _10067_ _10066_ _10065_ VGND VGND VPWR VPWR _10069_ sky130_fd_sc_hd__and3_1
XFILLER_145_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18126_ _09242_ _08970_ net605 _08969_ net779 VGND VGND VPWR VPWR _08974_ sky130_fd_sc_hd__o2111ai_4
X_15338_ _06095_ _06229_ _06230_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_117_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18057_ net615 net774 VGND VGND VPWR VPWR _08906_ sky130_fd_sc_hd__nand2_1
X_15269_ net739 a_h\[15\] VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__nand2_1
X_17008_ _07722_ net144 _07718_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__o21ai_1
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18959_ _09708_ _09634_ _09707_ VGND VGND VPWR VPWR _09851_ sky130_fd_sc_hd__a21boi_4
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer12 b_l\[4\] VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer45 net841 VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer34 _08777_ VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer23 net819 VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__buf_2
Xrebuffer78 net874 VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer56 _03953_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer67 net861 VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer89 net611 VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20783_ clknet_leaf_26_clk _00423_ VGND VGND VPWR VPWR a_l\[5\] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer102 a_l\[11\] VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_50_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer113 net909 VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer135 net684 VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__buf_4
Xrebuffer146 net942 VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer124 b_l\[0\] VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer157 _04409_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__buf_4
XFILLER_2_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold550 term_high\[55\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 term_high\[58\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap280 _07128_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__buf_6
XFILLER_116_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold572 _01257_ VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap291 net292 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20217_ net727 net548 VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__nand2_1
XFILLER_131_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20148_ _01316_ _01384_ _01382_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__nand3_1
XFILLER_106_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12970_ _02502_ _02589_ net659 net478 _03895_ VGND VGND VPWR VPWR _03897_ sky130_fd_sc_hd__o2111ai_1
X_20079_ _01292_ _01306_ _01308_ VGND VGND VPWR VPWR _01313_ sky130_fd_sc_hd__nand3b_1
XFILLER_18_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11921_ _02851_ _02852_ _02854_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__nand3_1
X_11852_ _02762_ _02786_ _02787_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__nand3b_4
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14640_ _09384_ _09406_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_103_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _01821_ _01824_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _05469_ _05470_ _09362_ _09406_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__o2bb2a_1
X_16310_ _07060_ _07181_ _07182_ net797 VGND VGND VPWR VPWR _07185_ sky130_fd_sc_hd__a31o_1
X_11783_ _02624_ _02638_ _02622_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__a21oi_2
X_13522_ _04429_ _04409_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_52_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_14_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17290_ _08152_ _08153_ _08155_ _08010_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__o2bb2ai_1
X_10734_ net467 _01763_ _01764_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_136_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16241_ net950 net515 _07112_ _07114_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__a22o_1
X_10665_ _01703_ _01704_ _01705_ _01700_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__a2bb2o_1
X_13453_ _04362_ _04363_ _04335_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__a21oi_2
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16172_ _07047_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__inv_2
X_12404_ _03331_ _03332_ _03333_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__a21o_1
X_13384_ _04294_ _04295_ VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__nand2_1
XFILLER_126_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10596_ _09690_ net1193 VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__and2_1
X_12335_ _03256_ _03266_ _03267_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__nand3_2
X_15123_ net733 net651 VGND VGND VPWR VPWR _06020_ sky130_fd_sc_hd__nand2_1
XFILLER_142_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12266_ _03196_ net398 VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__nand2_1
X_19931_ _01108_ _01146_ _01147_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__nand3_2
X_15054_ _05933_ _05935_ _05937_ _05949_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__o211ai_2
X_11217_ net681 net519 VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__nand2_2
X_12197_ net653 net508 VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__nand2_2
Xoutput70 net70 VGND VGND VPWR VPWR p[13] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19862_ _01075_ _01076_ _01077_ VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__a21o_1
X_14005_ _04888_ _04904_ _04906_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__nand3_1
Xoutput92 net92 VGND VGND VPWR VPWR p[33] sky130_fd_sc_hd__buf_2
X_11148_ net465 _02089_ _02076_ _02087_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__o211ai_2
X_18813_ _09676_ _09677_ net299 _09700_ VGND VGND VPWR VPWR _09706_ sky130_fd_sc_hd__o2bb2ai_1
Xoutput81 net81 VGND VGND VPWR VPWR p[23] sky130_fd_sc_hd__buf_2
X_19793_ net589 net725 VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_147_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15956_ _06719_ _06740_ _06827_ _06828_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__a2bb2oi_1
X_11079_ net697 net691 net1109 net519 VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__nand4_2
X_18744_ _09626_ _09627_ _09628_ VGND VGND VPWR VPWR _09631_ sky130_fd_sc_hd__a21o_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15887_ _09253_ _09581_ _06760_ _06762_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__o211ai_4
X_18675_ _09410_ _09411_ net737 _09217_ _09553_ VGND VGND VPWR VPWR _09556_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_19_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14907_ _05802_ _05804_ _05675_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__nand3_2
X_17626_ net560 net494 VGND VGND VPWR VPWR _08490_ sky130_fd_sc_hd__nand2_1
X_14838_ _05728_ _05734_ _05736_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__o21ai_2
XFILLER_24_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17557_ _08413_ _08415_ _08418_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_43_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_8
X_14769_ _05596_ _05636_ _05638_ _05597_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__a31oi_4
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16508_ net1004 net541 _07376_ _07378_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__a22o_1
X_17488_ _08336_ _08340_ _08351_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__o21ai_1
X_16439_ _07266_ _07267_ _07269_ _07270_ _07258_ VGND VGND VPWR VPWR _07312_ sky130_fd_sc_hd__a32o_2
X_19227_ _09874_ _09877_ _09900_ _10123_ VGND VGND VPWR VPWR _10125_ sky130_fd_sc_hd__o211ai_2
XFILLER_9_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19158_ _10041_ _10044_ _10045_ VGND VGND VPWR VPWR _10051_ sky130_fd_sc_hd__and3_1
XFILLER_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18109_ net458 _06401_ _08956_ VGND VGND VPWR VPWR _08957_ sky130_fd_sc_hd__a21o_1
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19089_ _05044_ _06441_ net411 _09766_ _09768_ VGND VGND VPWR VPWR _09980_ sky130_fd_sc_hd__o2111a_1
XFILLER_132_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_99_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20002_ _09340_ _01111_ _01109_ _01113_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__o22ai_2
XFILLER_143_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_34_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_146_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20766_ clknet_leaf_59_clk _00406_ VGND VGND VPWR VPWR a_h\[4\] sky130_fd_sc_hd__dfxtp_4
X_10450_ term_mid\[43\] term_high\[43\] _01613_ _01614_ VGND VGND VPWR VPWR _01615_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_118_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ clknet_leaf_4_clk _00337_ VGND VGND VPWR VPWR p_hl\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_10_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10381_ term_mid\[34\] term_high\[34\] VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__xor2_2
XTAP_TAPCELL_ROW_131_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12120_ net682 net679 net499 net492 VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__nand4_2
Xhold380 p_hh_pipe\[5\] VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12051_ _02984_ _02972_ _02983_ VGND VGND VPWR VPWR _02986_ sky130_fd_sc_hd__nand3_2
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11002_ net702 net697 net1109 net519 VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__nand4_2
Xhold391 p_ll_pipe\[1\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15810_ _06688_ _06675_ _06687_ VGND VGND VPWR VPWR _06689_ sky130_fd_sc_hd__nand3_2
X_16790_ _07655_ net344 _07636_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__a21oi_2
XFILLER_133_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15741_ net1110 _06595_ _06614_ _06616_ VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__o211ai_2
X_12953_ net659 net1015 net463 _03814_ VGND VGND VPWR VPWR _03880_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_5_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _02772_ _02836_ net692 net489 _02835_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o2111ai_2
X_15672_ _06550_ _06551_ _06513_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__nand3_2
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18460_ _09315_ _09320_ _09321_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__o21a_1
X_17411_ _08022_ _08159_ _08026_ _07879_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__nand4_1
X_12884_ _03810_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__nand2_1
X_14623_ _05385_ net709 b_l\[15\] VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_25_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
X_11835_ net687 net497 VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__nand2_2
X_18391_ _09244_ _09245_ _09232_ VGND VGND VPWR VPWR _09246_ sky130_fd_sc_hd__and3_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11766_ _02626_ _02630_ net462 VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__a21oi_1
X_17342_ net554 net969 VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__and2_1
XFILLER_13_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14554_ net1000 _05291_ _05452_ _05453_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__nand4_2
X_17273_ _08138_ _08139_ _08040_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__nand3_1
X_10717_ _01747_ _01749_ _01750_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__o21ba_1
X_13505_ net785 net673 net666 net1058 VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__a22o_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14485_ b_l\[15\] net709 _05383_ _05385_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__a22oi_2
X_11697_ net462 _02629_ net1048 net518 VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o211ai_1
X_16224_ _07096_ _07097_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__nand2_2
X_13436_ _04283_ _04288_ _04285_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__a21oi_1
X_19012_ _09747_ _09761_ VGND VGND VPWR VPWR _09903_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_24_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer3 net798 VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__clkbuf_2
X_10648_ p_hl\[4\] p_lh\[4\] VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__and2_1
X_10579_ net793 net1224 VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__and2_1
X_16155_ _09624_ _09635_ _06402_ _07029_ _07030_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__o32a_4
X_13367_ _04272_ _04274_ _04271_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12318_ _03249_ _03250_ _03251_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__o21a_1
X_16086_ net613 net607 net512 net505 VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__nand4_2
X_13298_ _04210_ _04209_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__nand2_1
X_15106_ _05910_ _05907_ _05999_ _06001_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__a211oi_4
X_12249_ _02833_ _03054_ _03050_ _03052_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_71_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19914_ net332 _01124_ _01130_ _01131_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__o2bb2ai_1
X_15037_ _05824_ _05923_ _05929_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__o2bb2ai_1
XTAP_TAPCELL_ROW_71_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19845_ _01059_ _01060_ _09231_ _09384_ VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__o2bb2ai_2
X_16988_ _07857_ net472 net843 _07856_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__nand4_1
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19776_ _00983_ _00984_ _09264_ _09340_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__o2bb2ai_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15939_ _06784_ net283 VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__nand2_1
X_18727_ net447 _09611_ _09600_ _09610_ VGND VGND VPWR VPWR _09612_ sky130_fd_sc_hd__o211ai_2
XFILLER_37_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18658_ _09534_ _09535_ VGND VGND VPWR VPWR _09538_ sky130_fd_sc_hd__nand2_2
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
X_17609_ _08413_ _08467_ _08468_ net414 VGND VGND VPWR VPWR _08473_ sky130_fd_sc_hd__a31o_1
X_18589_ _09359_ _09448_ _09459_ _09461_ VGND VGND VPWR VPWR _09462_ sky130_fd_sc_hd__o211ai_4
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20620_ clknet_leaf_42_clk _00260_ VGND VGND VPWR VPWR p_ll_pipe\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_138_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_82_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20551_ clknet_leaf_54_clk _00191_ VGND VGND VPWR VPWR mid_sum\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_146_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20482_ clknet_leaf_43_clk _00122_ VGND VGND VPWR VPWR term_mid\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_133_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11620_ _02348_ _02350_ _02553_ _02554_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__o211ai_1
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11551_ _02483_ _02485_ _02482_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_41_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10502_ term_high\[52\] term_high\[53\] term_high\[54\] VGND VGND VPWR VPWR _01657_
+ sky130_fd_sc_hd__and3_1
X_20749_ clknet_leaf_44_clk _00389_ VGND VGND VPWR VPWR p_ll\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11482_ _02270_ _02309_ _02310_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_21_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _05153_ _05154_ _05170_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__o21ai_4
X_10433_ _01597_ _01598_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__o21a_1
X_13221_ net784 net710 net704 net787 VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__a22o_1
Xwire568 net569 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__buf_12
XFILLER_109_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13152_ _09515_ _09679_ _04072_ net320 VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__o22a_1
XFILLER_6_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10364_ _01354_ _01364_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__nor2_1
XFILLER_128_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12103_ net358 _02875_ _02873_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__a21bo_1
XFILLER_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17960_ net623 net627 _04133_ VGND VGND VPWR VPWR _08813_ sky130_fd_sc_hd__and3_1
X_13083_ _03964_ _03904_ _04007_ _04005_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o2bb2ai_2
X_10295_ term_low\[21\] term_mid\[21\] VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__nand2_1
X_12034_ _02916_ _02880_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__nand2_2
X_17891_ net874 net938 net484 net480 _08720_ VGND VGND VPWR VPWR _08750_ sky130_fd_sc_hd__a41o_1
X_16911_ net571 net513 VGND VGND VPWR VPWR _07781_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_53_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16842_ _07710_ _07711_ _07703_ _07704_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__o211ai_2
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19630_ _00780_ _00828_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_144_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19561_ _00653_ _00744_ _00743_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_144_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16773_ _07641_ _07642_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__nand2_2
X_18512_ _09374_ _09375_ _09155_ _09275_ VGND VGND VPWR VPWR _09378_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13985_ net778 net656 VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__and2_1
X_15724_ _06601_ _06602_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__nand2_2
X_12936_ _03804_ _03805_ _03857_ net175 VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__nand4_1
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ net274 _00484_ _00452_ _00675_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__nand4_4
X_15655_ net624 net522 VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__nand2_1
X_12867_ _03795_ _03794_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__and2_1
X_18443_ _09298_ _09225_ _09214_ _09185_ VGND VGND VPWR VPWR _09303_ sky130_fd_sc_hd__a22oi_1
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11818_ _02752_ _02753_ _02719_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__a21oi_1
X_15586_ net628 net607 net1041 net522 VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__and4_1
X_18374_ _09131_ _09171_ _09169_ VGND VGND VPWR VPWR _09227_ sky130_fd_sc_hd__a21oi_2
XFILLER_61_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14606_ _05506_ _05507_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__nand2_1
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17325_ _08187_ _08189_ _08191_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__a21oi_4
X_12798_ _03528_ _03679_ _03665_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__o22ai_2
X_14537_ _04988_ net636 net778 VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__and3_1
X_11749_ _02684_ _02685_ _02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__nand3_1
XFILLER_147_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17256_ _08093_ _08118_ _08120_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__nand3_4
X_14468_ _05361_ _05369_ _05367_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__o21ai_1
X_16207_ _09166_ _09657_ _07074_ _07076_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__o211ai_2
X_17187_ net559 net509 VGND VGND VPWR VPWR _08055_ sky130_fd_sc_hd__nand2_2
X_13419_ _04327_ _04261_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__nand2_1
X_14399_ net756 net662 VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__nand2_1
XFILLER_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16138_ _06977_ _07011_ _07013_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__nand3_4
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16069_ _06937_ _06938_ _06942_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__nand3_1
XFILLER_103_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_5_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_57_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19828_ _01039_ _01037_ _01036_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__nand3b_4
Xclone8 net1020 net772 VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__nand2_8
X_19759_ _00858_ _00965_ _00966_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__nand3_4
XFILLER_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20603_ clknet_leaf_35_clk _00243_ VGND VGND VPWR VPWR p_ll_pipe\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20534_ clknet_leaf_47_clk _00174_ VGND VGND VPWR VPWR term_low\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20465_ clknet_leaf_14_clk _00105_ VGND VGND VPWR VPWR term_high\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_137_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20396_ clknet_leaf_47_clk _00036_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_126_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10982_ _01923_ net404 _01915_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__nand3_4
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13770_ _04675_ _04676_ _04655_ _04660_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__o211ai_2
X_12721_ _03646_ _03647_ _03650_ VGND VGND VPWR VPWR _03651_ sky130_fd_sc_hd__and3_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _03580_ _03416_ _03412_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__nand3b_2
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ _06292_ _06296_ _06329_ _06330_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__a22o_1
X_11603_ _02536_ _02538_ _02519_ _02521_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__o211ai_1
XFILLER_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12583_ _03151_ _03420_ _03511_ _03512_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a2bb2oi_1
X_15371_ net722 net640 VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__nand2_1
X_11534_ _02467_ _02469_ _02347_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__o21bai_4
X_17110_ _07963_ _07964_ _07974_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__nand3_1
X_18090_ _08935_ _08938_ _08899_ VGND VGND VPWR VPWR _08939_ sky130_fd_sc_hd__a21oi_1
Xwire321 _03524_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__buf_1
X_14322_ _05050_ _05065_ _05063_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__o21a_1
X_11465_ _09406_ _09613_ _02403_ _02404_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__o211ai_2
X_17041_ net418 _07904_ _07905_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__nand3_1
Xwire354 _03439_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_6
Xwire365 _00180_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14253_ _04982_ _04989_ _04985_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__a21oi_1
X_10416_ _01579_ _01583_ _01585_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__o21ai_1
XFILLER_137_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire398 _03180_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_1
X_13204_ _04111_ _04087_ _04109_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__or3b_1
X_11396_ _02251_ _02311_ _02312_ _02315_ _02249_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__a32oi_4
X_14184_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__inv_2
XFILLER_140_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13135_ _04019_ _04058_ _04022_ _04057_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__nand4_1
X_10347_ term_low\[29\] term_mid\[29\] VGND VGND VPWR VPWR _01192_ sky130_fd_sc_hd__and2_1
X_18992_ net598 net1091 VGND VGND VPWR VPWR _09883_ sky130_fd_sc_hd__nand2_2
XFILLER_140_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17943_ net170 VGND VGND VPWR VPWR _08800_ sky130_fd_sc_hd__inv_2
X_13066_ _03940_ _03943_ _03938_ VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__o21ai_1
X_10278_ _10158_ _10115_ net797 VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__a21oi_1
X_12017_ _02950_ _02951_ _02821_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__and3_1
X_17874_ _08728_ _08729_ _08733_ VGND VGND VPWR VPWR _08734_ sky130_fd_sc_hd__o21ai_2
Xclone222 net1028 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__clkbuf_16
X_19613_ _00808_ _00811_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__nand2_1
Xclone266 net544 VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__clkbuf_16
Xclone255 net1059 VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__clkbuf_16
X_16825_ _07545_ _07548_ _07691_ _07692_ VGND VGND VPWR VPWR _07696_ sky130_fd_sc_hd__o211ai_4
Xclone244 net543 VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__clkbuf_16
X_16756_ _07620_ _07621_ _07623_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__nand3_2
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19544_ _00734_ _00736_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__nor2_1
X_13968_ net762 net670 VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__nand2_1
X_15707_ net624 net515 VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__nand2_1
XFILLER_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12919_ _03844_ _03845_ _03808_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a21oi_1
X_19475_ _00458_ net579 b_l\[8\] VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__and3_1
X_16687_ _07555_ _07557_ _07489_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__a21o_1
X_18426_ _09282_ _09283_ _09267_ VGND VGND VPWR VPWR _09284_ sky130_fd_sc_hd__a21oi_1
X_13899_ _04800_ _04802_ _04774_ _04776_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__o211ai_2
X_15638_ net616 net527 VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_14_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15569_ _06447_ _06449_ _06435_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__a21oi_1
X_18357_ _09020_ _09096_ net149 _09208_ VGND VGND VPWR VPWR _09209_ sky130_fd_sc_hd__o31a_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17308_ net449 _08170_ _08168_ VGND VGND VPWR VPWR _08175_ sky130_fd_sc_hd__o21bai_2
X_18288_ net610 net764 VGND VGND VPWR VPWR _09134_ sky130_fd_sc_hd__nand2_1
XFILLER_119_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17239_ net573 net498 net493 net582 VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__a22oi_2
Xmax_cap621 net622 VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__buf_12
Xmax_cap632 a_l\[0\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_8
Xmax_cap654 a_h\[11\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__buf_12
Xmax_cap643 net907 VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__buf_8
X_20250_ _01490_ _01449_ _01448_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_110_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap665 net669 VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__buf_12
Xmax_cap676 net677 VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__buf_8
X_20181_ _01367_ _01374_ _01377_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_23_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap698 a_h\[3\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__buf_6
XFILLER_103_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_32_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20517_ clknet_leaf_41_clk _00157_ VGND VGND VPWR VPWR term_low\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_107_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20448_ clknet_leaf_18_clk _00088_ VGND VGND VPWR VPWR term_high\[40\] sky130_fd_sc_hd__dfxtp_1
X_11250_ _02107_ _02190_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__nand2_1
XFILLER_107_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_134_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11181_ _02035_ net363 _02033_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__a21o_1
X_20379_ clknet_leaf_32_clk _00019_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfxtp_1
XFILLER_79_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10201_ net548 VGND VGND VPWR VPWR _09373_ sky130_fd_sc_hd__inv_6
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14940_ net726 net723 net677 net861 VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__nand4_2
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14871_ _05769_ _05770_ _05667_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_141_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ _07470_ _07478_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__nand2_1
X_17590_ _08448_ _08450_ _08373_ VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__nand3_1
X_13822_ _04617_ _04604_ _04599_ _04605_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_16_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16541_ _07413_ _07412_ _07350_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__a21oi_2
X_13753_ net714 net731 VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__nand2_1
X_10965_ net707 net702 net1109 net1052 VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_106_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12704_ _03631_ _03633_ VGND VGND VPWR VPWR _03634_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16472_ _07338_ _07339_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__nand2_1
X_13684_ net777 net666 VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__nand2_2
X_10896_ net794 net1174 VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__and2_1
X_19260_ _10039_ _10049_ _10052_ VGND VGND VPWR VPWR _10161_ sky130_fd_sc_hd__nand3_2
XFILLER_129_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12635_ _03395_ _03407_ VGND VGND VPWR VPWR _03566_ sky130_fd_sc_hd__nand2_2
X_18211_ _09049_ _09055_ _09054_ VGND VGND VPWR VPWR _09058_ sky130_fd_sc_hd__o21ai_2
X_19191_ net598 net738 VGND VGND VPWR VPWR _10087_ sky130_fd_sc_hd__nand2_1
X_15423_ _06095_ _06229_ _06272_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_139_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _03497_ _03495_ net65 VGND VGND VPWR VPWR _03498_ sky130_fd_sc_hd__a21oi_1
X_18142_ _08986_ net764 net623 VGND VGND VPWR VPWR _08990_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_61_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _06244_ _06246_ _06241_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__nand3_2
XFILLER_12_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11517_ _02453_ _02454_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__nand2_2
XFILLER_8_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14305_ _05053_ _05207_ b_l\[11\] net695 _05206_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__o2111ai_4
XFILLER_11_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18073_ _08920_ _08921_ net779 net611 VGND VGND VPWR VPWR _08922_ sky130_fd_sc_hd__and4_1
X_12497_ net906 b_h\[8\] VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__nand2_1
X_15285_ _06153_ _06155_ _06175_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11448_ net360 _02288_ _02289_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__a21boi_1
X_17024_ _09188_ _09679_ _07890_ _07891_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__o22ai_2
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14236_ _05134_ _05136_ _05120_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__a21o_1
X_11379_ _02249_ _02315_ _02316_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__nand3_2
X_14167_ _05070_ _05064_ _05041_ _05071_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__o211a_1
X_13118_ net641 net634 net1151 net999 VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__nand4_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18975_ _09852_ _09739_ VGND VGND VPWR VPWR _09866_ sky130_fd_sc_hd__nand2_1
X_14098_ _04998_ _04979_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__nand2_1
X_17926_ _08782_ _08783_ _08758_ VGND VGND VPWR VPWR _08784_ sky130_fd_sc_hd__a21oi_1
X_13049_ _03958_ _03972_ _03973_ VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__nand3_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17857_ _08712_ _08715_ _08717_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__o21a_1
XFILLER_27_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16808_ _07666_ _07673_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__nand2_1
XFILLER_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17788_ _08580_ _08583_ _08587_ VGND VGND VPWR VPWR _08650_ sky130_fd_sc_hd__o21ai_1
X_19527_ _00586_ _00587_ _00685_ _00694_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__o22ai_1
X_16739_ _09210_ _09646_ _07609_ VGND VGND VPWR VPWR _07610_ sky130_fd_sc_hd__o21ai_1
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19458_ _10177_ _00642_ _10036_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__nand3_4
XFILLER_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18409_ _09229_ _09262_ _09263_ VGND VGND VPWR VPWR _09266_ sky130_fd_sc_hd__nand3_4
XFILLER_50_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19389_ _10156_ _00565_ _00566_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__nand3_2
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer317 _07035_ VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer306 net236 VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__buf_1
Xrebuffer328 _04259_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__buf_2
XFILLER_135_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20302_ _01546_ net152 VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__nor2_1
Xmax_cap462 _02627_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__buf_4
Xmax_cap451 _07967_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_2
X_20233_ _01474_ _01476_ _01468_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__o21ai_1
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap484 net486 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_12
Xmax_cap495 b_h\[10\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__buf_12
Xmax_cap473 net474 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_6
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_89_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20164_ _01402_ _01403_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__nand2_1
X_20095_ _09275_ _09384_ _01326_ _01327_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__o211ai_2
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10750_ p_hl\[20\] p_lh\[20\] VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_36_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10681_ p_hl\[9\] p_lh\[9\] VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__xnor2_1
X_12420_ _03350_ _03351_ a_h\[3\] net474 VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__nand4_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12351_ _03280_ _03282_ _03278_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__a21oi_2
X_11302_ net712 net983 net975 net491 VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__and4_2
X_12282_ _03169_ _03171_ _03206_ _03208_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__nand4_1
XFILLER_4_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15070_ _05819_ _05903_ _05965_ _05966_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_134_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11233_ net1061 net1024 _02169_ _02171_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__a22o_1
XFILLER_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021_ _04707_ _04923_ _04925_ _04708_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_20_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_122_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11164_ net706 net507 VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__nand2_1
X_15972_ net496 net491 net849 _06848_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__a31o_1
X_11095_ net707 net1018 net507 net712 VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__a22oi_1
XFILLER_95_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18760_ net775 net1146 net581 net576 _09639_ VGND VGND VPWR VPWR _09649_ sky130_fd_sc_hd__a41o_1
X_17711_ _08569_ _08572_ _08573_ VGND VGND VPWR VPWR _08574_ sky130_fd_sc_hd__a21oi_1
X_18691_ _09566_ _09571_ _09567_ VGND VGND VPWR VPWR _09574_ sky130_fd_sc_hd__nand3_2
X_14923_ net739 net655 VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__nand2_1
XFILLER_75_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17642_ _08501_ _08503_ _08488_ VGND VGND VPWR VPWR _08506_ sky130_fd_sc_hd__o21bai_1
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14854_ net285 _05633_ _05753_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__nand3_4
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11997_ _02932_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__inv_2
X_17573_ _08436_ _08437_ _08432_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__a21oi_1
XFILLER_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14785_ net756 net750 net649 net642 VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__nand4_2
X_13805_ _09264_ _09417_ _04632_ _04707_ _04711_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__o221ai_2
X_10948_ _01892_ _01893_ _01894_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__a21oi_2
X_16524_ _07391_ _07393_ net583 net516 VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__o211a_1
X_13736_ net393 _04642_ _04628_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__a21o_1
X_19312_ _10032_ _10058_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__nand2_1
X_16455_ _09624_ _07325_ net1032 net620 _07324_ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__o2111ai_4
X_19243_ _09981_ net717 net630 _09978_ VGND VGND VPWR VPWR _10143_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_14_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10879_ net794 net1162 VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__and2_1
X_13667_ _04391_ _04392_ _04571_ _04573_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__o211ai_2
X_15406_ _06254_ _06257_ _06297_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_14_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16386_ a_l\[7\] net513 VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__nand2_1
X_12618_ _03542_ _03543_ net436 VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__nand3_2
X_13598_ net772 net675 VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__nand2_1
X_19174_ _09924_ _09959_ _09957_ VGND VGND VPWR VPWR _10068_ sky130_fd_sc_hd__a21oi_4
XFILLER_129_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12549_ _03347_ _03354_ VGND VGND VPWR VPWR _03481_ sky130_fd_sc_hd__nand2_1
X_18125_ _08969_ _08971_ _08965_ VGND VGND VPWR VPWR _08973_ sky130_fd_sc_hd__a21bo_1
X_15337_ _06095_ _06229_ _06230_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__o21a_1
XFILLER_8_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_1 _00051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18056_ net623 net769 VGND VGND VPWR VPWR _08905_ sky130_fd_sc_hd__nand2_1
X_15268_ net739 net733 net641 a_h\[15\] VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__nand4_4
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_144_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17007_ _07589_ _07713_ _07714_ _07723_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__a31oi_1
X_14219_ net750 net670 VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__nand2_1
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15199_ net733 net913 VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_74_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18958_ _09848_ _09849_ VGND VGND VPWR VPWR _09850_ sky130_fd_sc_hd__nand2_1
X_17909_ _08767_ VGND VGND VPWR VPWR _08768_ sky130_fd_sc_hd__inv_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18889_ _09779_ _09780_ _09776_ VGND VGND VPWR VPWR _09781_ sky130_fd_sc_hd__a21o_1
Xrebuffer46 a_l\[2\] VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_67_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer35 _09851_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer13 b_l\[4\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer24 net820 VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer79 net874 VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer57 net648 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer68 net861 VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20782_ clknet_leaf_19_clk _00422_ VGND VGND VPWR VPWR a_l\[4\] sky130_fd_sc_hd__dfxtp_4
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer103 net899 VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer136 net932 VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer114 net909 VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer158 _06624_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__buf_2
XFILLER_123_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold551 p_ll\[30\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 p_ll\[27\] VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap270 _01243_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__buf_1
Xmax_cap281 net282 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__buf_1
XFILLER_104_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap292 _03451_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_2
X_20216_ _01218_ _01361_ _01419_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__o21ai_1
Xhold573 term_mid\[26\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20147_ _01316_ _01384_ _01382_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__and3_1
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20078_ _01287_ _01290_ _01305_ net331 VGND VGND VPWR VPWR _01312_ sky130_fd_sc_hd__o22ai_2
X_11920_ _02852_ _02854_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__nand2_1
XFILLER_85_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11851_ _02785_ _02762_ _02784_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__nand3_1
X_11782_ _02717_ _02718_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_103_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _01816_ _01822_ _01823_ _01814_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__o22ai_1
XFILLER_82_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _05330_ _05466_ net720 net699 _05470_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__o2111ai_4
XFILLER_26_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10733_ _01763_ net467 net796 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a21oi_1
X_13521_ _04427_ _04428_ _04409_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_45_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16240_ net950 net515 _07112_ _07114_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__a22oi_1
X_10664_ p_hl\[5\] p_lh\[5\] _01705_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__o21ai_1
X_13452_ _04359_ _04345_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nand2_1
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16171_ _07046_ net260 _07044_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__nand3_2
X_10595_ _09690_ net1188 VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__and2_1
X_12403_ _03331_ _03332_ _03333_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a21oi_1
X_13383_ _04292_ _04281_ _04291_ VGND VGND VPWR VPWR _04295_ sky130_fd_sc_hd__nand3_2
X_12334_ _03260_ _03263_ _03257_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__a21o_1
X_15122_ net739 net909 VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__nand2_2
XFILLER_126_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19930_ _01108_ _01148_ _01151_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__nand3b_2
X_15053_ _05945_ _05947_ _05938_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12265_ _03181_ _03194_ _03195_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nand3_1
XFILLER_99_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14004_ _04880_ _04881_ _04903_ _04905_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__o22ai_2
X_11216_ _02067_ _02156_ VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__nand2_2
X_12196_ _02978_ _03128_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__nand2_2
X_19861_ _01075_ _01076_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__a21oi_2
Xoutput93 net93 VGND VGND VPWR VPWR p[34] sky130_fd_sc_hd__buf_2
X_11147_ _02005_ _02075_ net465 _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__o2bb2ai_2
Xoutput71 net71 VGND VGND VPWR VPWR p[14] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18812_ net1031 net1081 _09698_ _09701_ VGND VGND VPWR VPWR _09705_ sky130_fd_sc_hd__nand4_2
X_19792_ _00883_ _01002_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__nand2_1
Xoutput82 net82 VGND VGND VPWR VPWR p[24] sky130_fd_sc_hd__buf_2
X_18743_ _09626_ _09627_ _09628_ VGND VGND VPWR VPWR _09630_ sky130_fd_sc_hd__nand3_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15955_ _06832_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__inv_2
X_11078_ _01945_ _02020_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__nand2_1
X_15886_ _06760_ _06762_ _09253_ _09581_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_91_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18674_ _09545_ _09549_ _09551_ _09547_ VGND VGND VPWR VPWR _09555_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_19_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14906_ _05801_ _05803_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__nor2_1
X_17625_ _08309_ _08395_ _08394_ VGND VGND VPWR VPWR _08489_ sky130_fd_sc_hd__a21oi_1
XFILLER_63_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14837_ _05736_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__inv_2
X_17556_ _08313_ _08326_ _08413_ _08415_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__nand4_1
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16507_ _07376_ _07378_ _09340_ _09581_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__o2bb2a_1
X_14768_ _05596_ _05636_ _05638_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__nand3_1
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17487_ _08336_ _08340_ _08351_ _08350_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__a2bb2o_2
X_13719_ _09406_ _09417_ _04260_ _04492_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__o31a_2
X_14699_ _05417_ net1060 _05425_ _05428_ _05432_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__a32oi_4
X_16438_ _06961_ _07129_ _07133_ _07272_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__o211a_1
X_19226_ _09874_ _09877_ _09900_ _10123_ VGND VGND VPWR VPWR _10124_ sky130_fd_sc_hd__o211a_1
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16369_ net559 net544 net523 net583 VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__a22o_1
X_19157_ _10045_ _10044_ _10041_ VGND VGND VPWR VPWR _10049_ sky130_fd_sc_hd__a21o_1
X_18108_ net626 net759 net754 net630 VGND VGND VPWR VPWR _08956_ sky130_fd_sc_hd__a22oi_1
XFILLER_118_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19088_ _09744_ net411 _09766_ _09768_ VGND VGND VPWR VPWR _09979_ sky130_fd_sc_hd__a22o_1
X_18039_ _08886_ _08887_ _08831_ VGND VGND VPWR VPWR _08889_ sky130_fd_sc_hd__nand3_1
X_20001_ _01110_ _01218_ _01216_ _01223_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__o211ai_1
XFILLER_100_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20765_ clknet_leaf_1_clk _00405_ VGND VGND VPWR VPWR a_h\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20696_ clknet_leaf_4_clk _00336_ VGND VGND VPWR VPWR p_hl\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10380_ _01513_ _01524_ _01534_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_131_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold370 p_ll\[6\] VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12050_ _02984_ _02972_ _02983_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__and3_1
Xhold381 p_ll\[9\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net697 net1109 VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__nand2_1
Xhold392 term_low\[1\] VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15740_ _06619_ VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__inv_2
XFILLER_93_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12952_ net944 net474 VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _02835_ _02837_ _09417_ _09646_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__o2bb2ai_1
X_15671_ _06482_ _06488_ _06512_ _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__o211ai_2
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17410_ _07584_ _08024_ _08274_ _07586_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__nand4_4
X_12883_ net654 b_h\[12\] VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__nand2_1
X_14622_ _05411_ _05519_ _05520_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__nand3_4
X_11834_ net692 net492 VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__nand2_1
X_18390_ _09155_ _09253_ net459 _07100_ _09238_ VGND VGND VPWR VPWR _09245_ sky130_fd_sc_hd__o221ai_4
XFILLER_60_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11765_ _02626_ _02630_ net462 VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__a21o_1
X_17341_ _08055_ _08207_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__nand2_2
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14553_ _05289_ _05438_ _05454_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__a21oi_2
X_11696_ net462 _02630_ net1048 net518 VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__and4b_1
X_17272_ _08138_ _08139_ _08040_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__and3_4
X_10716_ _01744_ _01748_ _01747_ net796 VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__a31o_1
X_13504_ net785 net673 net666 net1058 VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a22oi_1
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14484_ _05383_ _05385_ b_l\[15\] net709 VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__and4_1
XFILLER_146_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16223_ net572 net532 net528 net582 VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__a22oi_1
X_10647_ p_hl\[4\] p_lh\[4\] VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__nor2_1
X_13435_ _04283_ _04288_ _04285_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__a21o_1
X_19011_ _09605_ _09616_ _09755_ _09757_ _09747_ VGND VGND VPWR VPWR _09902_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_24_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer4 net800 VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd1_1
X_10578_ net793 net1307 VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__and2_1
X_16154_ _09166_ _09646_ _07027_ _07028_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__nor4_4
X_13366_ _09220_ _09395_ _01888_ net805 _04274_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_58_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12317_ _03250_ _03249_ net65 VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__a21oi_1
XFILLER_127_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16085_ net607 net505 VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__nand2_4
X_13297_ _04174_ _04178_ _04209_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__a21o_1
X_15105_ _05797_ _05906_ _05999_ _06001_ _05910_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__o221a_1
X_12248_ _03050_ net461 _03055_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__o21ai_1
X_19913_ _01130_ _01131_ VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__nor2_1
X_15036_ _05925_ _05928_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__nand2_1
XFILLER_123_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19844_ _00901_ _00907_ _00940_ _00946_ VGND VGND VPWR VPWR _01060_ sky130_fd_sc_hd__o211ai_2
X_12179_ _02954_ _02957_ _03110_ _03111_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__nand4_1
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16987_ _07621_ _07854_ _07853_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__a21o_1
XFILLER_84_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19775_ _00983_ _00984_ _09264_ _09340_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__o2bb2a_1
X_15938_ _06784_ _06787_ net283 VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__a21oi_1
XFILLER_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18726_ net619 net609 net743 net737 _09609_ VGND VGND VPWR VPWR _09611_ sky130_fd_sc_hd__a41o_1
X_18657_ net618 net743 net737 net621 VGND VGND VPWR VPWR _09536_ sky130_fd_sc_hd__a22oi_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15869_ _09166_ _09624_ _06744_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__o21a_1
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17608_ _09253_ _09679_ VGND VGND VPWR VPWR _08472_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18588_ net457 _06681_ _09451_ _09454_ VGND VGND VPWR VPWR _09461_ sky130_fd_sc_hd__o211ai_2
XFILLER_52_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17539_ _08397_ _08399_ _08394_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_82_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20550_ clknet_leaf_54_clk _00190_ VGND VGND VPWR VPWR mid_sum\[13\] sky130_fd_sc_hd__dfxtp_1
X_19209_ _10100_ _10075_ _10101_ VGND VGND VPWR VPWR _10106_ sky130_fd_sc_hd__nand3_4
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20481_ clknet_leaf_43_clk _00121_ VGND VGND VPWR VPWR term_mid\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_145_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11550_ _09449_ _09602_ _02486_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__o21ai_4
X_20748_ clknet_leaf_42_clk _00388_ VGND VGND VPWR VPWR p_ll\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10501_ net796 net1332 _01656_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__nor3_1
XFILLER_50_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ _02308_ _02307_ _02271_ _02310_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__a22oi_2
Xwire547 b_h\[0\] VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__buf_12
X_13220_ _01860_ _04134_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__or2_1
X_20679_ clknet_leaf_55_clk _00319_ VGND VGND VPWR VPWR p_hl\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10432_ _01595_ _01590_ _01589_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__a21oi_1
XFILLER_136_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13151_ _09515_ net320 _09679_ _04072_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__nor4_1
X_10363_ term_low\[31\] term_mid\[31\] VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__and2_1
X_12102_ _02971_ _03030_ _03032_ VGND VGND VPWR VPWR _03037_ sky130_fd_sc_hd__nand3_4
X_13082_ _04003_ _04004_ _04001_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12033_ _02937_ _02946_ _02933_ _02935_ VGND VGND VPWR VPWR _02968_ sky130_fd_sc_hd__o2bb2ai_1
X_16910_ net1069 net503 VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__nand2_1
XFILLER_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10294_ term_low\[21\] term_mid\[21\] VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__and2_1
XFILLER_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17890_ net796 _08748_ _08749_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__nor3_1
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16841_ _07710_ _07711_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_144_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16772_ net874 net534 net530 net558 VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__a22oi_4
XFILLER_93_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_69_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19560_ _09319_ _09340_ net457 _09297_ _09264_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__o32a_1
XFILLER_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_144_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ net607 net531 net527 net1090 VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__a22oi_1
XFILLER_92_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18511_ _09374_ _09375_ _09369_ VGND VGND VPWR VPWR _09377_ sky130_fd_sc_hd__a21o_1
X_13984_ _09155_ _09482_ _02502_ _04134_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__o22a_1
X_12935_ _03804_ _03805_ _03858_ VGND VGND VPWR VPWR _03863_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_29_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19491_ _00677_ _00678_ _00679_ net298 VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__a22oi_2
X_15654_ net628 net515 VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__nand2_2
X_12866_ _03790_ _03791_ _03793_ net793 VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__o31a_1
X_18442_ _09223_ _09224_ _09298_ VGND VGND VPWR VPWR _09302_ sky130_fd_sc_hd__o21ai_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15585_ net607 net521 VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__nand2_1
X_11817_ _02752_ _02753_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__nand2_1
X_18373_ _09126_ _09127_ _09170_ VGND VGND VPWR VPWR _09226_ sky130_fd_sc_hd__o21ai_1
X_14605_ _05505_ _05504_ _05413_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__nand3_4
X_17324_ _08061_ _08064_ _08063_ _08069_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__a22oi_4
X_12797_ _03670_ _03680_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__nand2_1
XFILLER_14_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14536_ _05280_ _05281_ net1000 VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__nand3_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11748_ _02554_ _02351_ _02552_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_78_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11679_ _02615_ _02607_ VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__nand2_1
X_17255_ _08122_ _08092_ _08121_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__nand3_4
X_14467_ _05362_ _05363_ _05219_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__and3_1
X_16206_ _07080_ _07064_ _07079_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__nand3_2
X_17186_ _07925_ _08052_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__nand2_4
X_13418_ net435 _04324_ _04325_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__nand3_1
X_14398_ net746 net670 VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__nand2_1
XFILLER_142_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16137_ _07005_ _07007_ _06990_ _06994_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__o211ai_2
XFILLER_115_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13349_ net714 net963 net1125 VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__and3_1
XFILLER_142_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16068_ _06745_ _06934_ _06936_ _06944_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__a31o_1
XFILLER_115_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_87_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15019_ _05812_ _05914_ _05813_ _05673_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__and4_1
XFILLER_96_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19827_ _00927_ _00937_ _01037_ _01036_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__a22o_1
XFILLER_110_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19758_ _00965_ _00966_ _00858_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18709_ _09588_ _09591_ _09593_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__a21boi_1
X_19689_ _00888_ _00889_ b_l\[5\] net548 VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__nand4_2
XFILLER_80_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20602_ clknet_leaf_35_clk _00242_ VGND VGND VPWR VPWR p_ll_pipe\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_96_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20533_ clknet_leaf_49_clk _00173_ VGND VGND VPWR VPWR term_low\[28\] sky130_fd_sc_hd__dfxtp_1
X_20464_ clknet_leaf_14_clk _00104_ VGND VGND VPWR VPWR term_high\[56\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_95_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20395_ clknet_leaf_36_clk _00035_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_87_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10981_ _01916_ _01925_ _01926_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__nand3_4
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12720_ _03541_ _03648_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__nand2_1
XFILLER_71_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12651_ _03411_ _03580_ _03581_ VGND VGND VPWR VPWR _03582_ sky130_fd_sc_hd__nand3_2
XFILLER_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11602_ _02519_ _02521_ _02540_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__a21o_1
XFILLER_90_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12582_ _09504_ _03510_ _03512_ VGND VGND VPWR VPWR _03513_ sky130_fd_sc_hd__o21ai_1
X_15370_ _06261_ _06262_ _06263_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11533_ _02468_ _02470_ _02243_ net402 VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__nand4_1
Xwire322 _03445_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_2
Xwire300 _09622_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_1
XFILLER_7_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire311 _05852_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__buf_1
X_14321_ _05223_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__nand2_1
X_11464_ _02395_ net507 net692 VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__nand3_1
X_17040_ _07900_ _07901_ _07903_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__nand3_1
Xwire366 _00986_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_1
X_14252_ _04982_ _04989_ _04985_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a21o_1
X_10415_ term_mid\[39\] term_high\[39\] VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__xor2_1
XFILLER_125_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13203_ _04087_ _04112_ VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__nor2_1
X_11395_ _02332_ net982 _02335_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__o21ba_1
X_14183_ _05087_ net431 net709 net724 VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__and4b_1
XFILLER_124_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_98_718 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13134_ _04055_ _04056_ _04049_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21o_1
X_18991_ net603 net738 VGND VGND VPWR VPWR _09882_ sky130_fd_sc_hd__nand2_2
X_10346_ _01106_ _01161_ _01172_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__a21oi_1
XFILLER_140_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17942_ _08797_ _08798_ VGND VGND VPWR VPWR _08799_ sky130_fd_sc_hd__xor2_1
X_13065_ _03988_ _03989_ _03957_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__a21bo_1
X_10277_ _10158_ _10115_ VGND VGND VPWR VPWR _10169_ sky130_fd_sc_hd__nand2_1
X_12016_ _02821_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__nand2_1
X_17873_ _08728_ _08729_ _08724_ VGND VGND VPWR VPWR _08733_ sky130_fd_sc_hd__a21oi_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16824_ _07693_ _07694_ _07629_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__a21oi_2
X_19612_ _00805_ _00807_ _00796_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__nand3_2
X_16755_ _07620_ _07621_ _07623_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__a21o_1
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclone267 net1066 VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__clkbuf_16
X_19543_ net765 net552 net548 net919 VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__a22oi_4
X_13967_ _04752_ _04754_ _04756_ _04741_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__a2bb2oi_2
X_16686_ _07550_ _07554_ _07557_ _07489_ VGND VGND VPWR VPWR _07558_ sky130_fd_sc_hd__o211ai_2
X_15706_ _06545_ net309 _06532_ _06530_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_73_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12918_ _03844_ _03845_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19474_ _00658_ _00657_ _00647_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__nand3_4
X_15637_ net607 net540 VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18425_ _09279_ _09280_ _09268_ VGND VGND VPWR VPWR _09283_ sky130_fd_sc_hd__nand3_2
X_13898_ _04797_ _04798_ _04668_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__a21oi_1
X_12849_ _03721_ _03724_ _03774_ _03776_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__o211ai_1
X_15568_ _06433_ _06434_ _06447_ _06449_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__o211ai_1
X_18356_ _09020_ _09096_ net149 _09207_ VGND VGND VPWR VPWR _09208_ sky130_fd_sc_hd__o22ai_4
X_18287_ net372 _09073_ _09074_ _09058_ VGND VGND VPWR VPWR _09133_ sky130_fd_sc_hd__a2bb2oi_2
X_17307_ _02338_ _07234_ _08168_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__o21ai_2
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14519_ _05419_ _05420_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nand2_2
X_15499_ net719 net716 net640 net635 _06387_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__a41o_1
XFILLER_147_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17238_ net573 net498 VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__nand2_1
Xmax_cap611 a_l\[4\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__buf_12
Xmax_cap600 net601 VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_6
X_17169_ _08035_ _08036_ _08032_ VGND VGND VPWR VPWR _08037_ sky130_fd_sc_hd__a21o_1
Xmax_cap622 net623 VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__buf_12
Xmax_cap644 net645 VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__buf_12
Xmax_cap633 net634 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__buf_8
XFILLER_131_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap688 a_h\[5\] VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__buf_12
Xmax_cap677 a_h\[7\] VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__buf_12
X_20180_ _01359_ _01363_ _01373_ _01376_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__o2bb2ai_1
Xmax_cap666 net667 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__buf_6
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap699 net701 VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_8
XFILLER_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20516_ clknet_leaf_41_clk _00156_ VGND VGND VPWR VPWR term_low\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_119_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20447_ clknet_leaf_27_clk _00087_ VGND VGND VPWR VPWR term_high\[39\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10200_ net720 VGND VGND VPWR VPWR _09362_ sky130_fd_sc_hd__clkinv_8
X_11180_ _02099_ _02101_ _02116_ _02118_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__nand4_1
X_20378_ clknet_leaf_33_clk _00018_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfxtp_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14870_ _05642_ _05646_ _05764_ _05765_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_141_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13821_ _04599_ _04605_ _04617_ _04604_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a2bb2oi_1
X_16540_ _07409_ _07367_ VGND VGND VPWR VPWR _07413_ sky130_fd_sc_hd__nand2_2
XFILLER_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13752_ _04586_ _04656_ _04658_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__nand3_4
XFILLER_16_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10964_ net707 net702 net1109 net1052 VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_106_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12703_ net680 net475 _03628_ _03629_ VGND VGND VPWR VPWR _03633_ sky130_fd_sc_hd__a22o_1
XFILLER_44_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16471_ _07338_ _07341_ _07339_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__a21o_1
X_18210_ _09049_ _09055_ _09054_ VGND VGND VPWR VPWR _09057_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13683_ net777 net666 VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__and2_1
X_10895_ net794 net1169 VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__and2_1
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12634_ _03535_ _03559_ _03561_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__nand3b_4
XFILLER_70_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19190_ net603 net732 VGND VGND VPWR VPWR _10086_ sky130_fd_sc_hd__nand2_2
X_15422_ _06312_ _06313_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_139_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _03372_ _03374_ _03370_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__o21ai_1
XFILLER_129_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18141_ net623 net764 _08986_ _08988_ VGND VGND VPWR VPWR _08989_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_61_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15353_ _09384_ _09482_ _06243_ _06245_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__o22ai_4
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11516_ net706 net698 net497 net492 VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__nand4_1
X_18072_ net790 net781 net605 net601 VGND VGND VPWR VPWR _08921_ sky130_fd_sc_hd__nand4_2
Xwire141 _01500_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
X_14304_ net740 net736 net690 net685 VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__nand4_2
XFILLER_12_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17023_ _02589_ _06605_ net377 _07770_ _07774_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__o2111ai_4
X_12496_ net653 b_h\[8\] VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__and2_1
X_15284_ _06172_ _06176_ _05999_ _06177_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__o211ai_2
Xwire163 _05649_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_6
Xwire152 _01547_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xwire174 _06054_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_1
X_11447_ _02282_ _02284_ _02287_ _02289_ _02302_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__a32oi_2
Xwire185 _09565_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
X_14235_ _05134_ _05136_ _05120_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__a21oi_2
X_11378_ _02316_ _02315_ _02249_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__a21o_1
XFILLER_125_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14166_ net350 _05066_ _05050_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__a21o_1
X_13117_ net641 net634 net1151 net999 VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__and4_1
X_10329_ term_low\[25\] term_mid\[25\] _00978_ _00870_ VGND VGND VPWR VPWR _00999_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18974_ _09861_ _09863_ VGND VGND VPWR VPWR _09865_ sky130_fd_sc_hd__nor2_1
X_14097_ _04974_ _04977_ _04978_ _04994_ _04997_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__o2111ai_1
X_17925_ a_l\[15\] net477 net473 net555 VGND VGND VPWR VPWR _08783_ sky130_fd_sc_hd__a22o_1
XFILLER_78_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13048_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__nand2_1
X_17856_ _08712_ _08715_ net796 VGND VGND VPWR VPWR _08717_ sky130_fd_sc_hd__a21oi_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16807_ _07666_ _07676_ _07677_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__nand3b_4
X_17787_ _08577_ _08585_ _08587_ VGND VGND VPWR VPWR _08649_ sky130_fd_sc_hd__o21bai_1
X_16738_ _02338_ _06761_ _07608_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__o21ai_1
X_14999_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__inv_2
X_19526_ _00580_ _00585_ _00584_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__a21oi_1
X_16669_ net379 _07536_ _07519_ _07538_ VGND VGND VPWR VPWR _07541_ sky130_fd_sc_hd__o211ai_4
X_19457_ _10036_ _10177_ _00640_ _00641_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__o2bb2ai_4
X_18408_ _09230_ _09260_ _09261_ VGND VGND VPWR VPWR _09265_ sky130_fd_sc_hd__nand3_4
X_19388_ _00567_ _10157_ _00568_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__nand3_4
XTAP_TAPCELL_ROW_17_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18339_ _09038_ _09042_ _09187_ VGND VGND VPWR VPWR _09190_ sky130_fd_sc_hd__a21oi_1
Xrebuffer318 b_h\[0\] VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer307 _08777_ VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__buf_1
Xrebuffer329 net1125 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_TAPCELL_ROW_79_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20301_ _01532_ _01536_ _01545_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__nor3b_1
XFILLER_146_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap452 _07752_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_92_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap463 _02588_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_6
X_20232_ _01472_ _01473_ _01469_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_92_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap485 net486 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_12
Xmax_cap474 b_h\[15\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_6
X_20163_ _01338_ _01342_ _01399_ _01400_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__nand4_1
XFILLER_131_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20094_ _01326_ _01327_ _01325_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__a21o_1
XFILLER_111_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10680_ _01710_ net469 _01715_ net797 _01718_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__a311oi_1
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12350_ _03278_ _03282_ _03280_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__and3_1
X_11301_ net983 net975 _09635_ _09177_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__o2bb2a_1
X_12281_ _03169_ _03171_ _03209_ _03211_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__nand4_2
XFILLER_5_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11232_ _02079_ _02170_ net1061 net1024 _02169_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o2111ai_4
X_14020_ net758 net752 net683 net676 VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__nand4_1
XFILLER_134_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11163_ _02037_ _02104_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__nand2_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15971_ net629 net496 _09635_ _09166_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__o2bb2a_1
X_11094_ net712 net707 net510 net507 VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__and4_1
XFILLER_121_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17710_ _08497_ _08492_ _08495_ VGND VGND VPWR VPWR _08573_ sky130_fd_sc_hd__o21ai_2
X_18690_ _09402_ _09567_ _09569_ VGND VGND VPWR VPWR _09573_ sky130_fd_sc_hd__nand3_4
X_14922_ net733 net663 VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__nand2_1
XFILLER_76_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17641_ _08488_ _08502_ _08504_ VGND VGND VPWR VPWR _08505_ sky130_fd_sc_hd__nand3_1
X_14853_ _05467_ _05604_ net389 VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__o21ai_2
XFILLER_76_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13804_ _04635_ _04708_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__nand2_2
X_11996_ _02855_ _02857_ _02925_ _02928_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__nand4_2
XFILLER_91_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17572_ _08301_ _08328_ _08331_ _08433_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__o211ai_4
XFILLER_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14784_ net756 net750 net649 net642 VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__and4_1
X_19311_ _00483_ _00485_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__nand2_2
X_10947_ _01868_ _01869_ _01872_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__o21ai_2
X_16523_ _07391_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__nor2_1
X_13735_ net393 _04642_ _04628_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16454_ net620 net487 VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__and2_1
X_13666_ _04393_ _04571_ _04573_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__nand3b_4
X_19242_ _10140_ _10141_ VGND VGND VPWR VPWR _10142_ sky130_fd_sc_hd__nand2_1
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10878_ _09690_ net1167 VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__and2_1
X_12617_ net436 _03545_ _03544_ VGND VGND VPWR VPWR _03548_ sky130_fd_sc_hd__nand3b_2
X_15405_ _06254_ _06257_ _06297_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__a21boi_1
X_19173_ _09924_ _09959_ _09956_ _09953_ VGND VGND VPWR VPWR _10067_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_TAPCELL_ROW_14_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _07258_ VGND VGND VPWR VPWR _07259_ sky130_fd_sc_hd__inv_2
X_18124_ net779 net605 _08969_ _08971_ VGND VGND VPWR VPWR _08972_ sky130_fd_sc_hd__a22oi_2
XPHY_EDGE_ROW_51_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13597_ net762 net689 VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__nand2_1
XFILLER_8_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12548_ _03463_ _03464_ _03476_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__nand3_2
X_15336_ _06162_ _06228_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__nand2_1
XFILLER_8_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_2 _00052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12479_ _03271_ _03409_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__nand3_2
X_18055_ net626 net764 VGND VGND VPWR VPWR _08904_ sky130_fd_sc_hd__nand2_1
X_15267_ net733 a_h\[15\] VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__nand2_1
XFILLER_144_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17006_ _07868_ _07869_ _07870_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__nand3_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14218_ net746 net676 VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__nand2_1
X_15198_ _06091_ _06092_ VGND VGND VPWR VPWR _06094_ sky130_fd_sc_hd__nand2_1
XFILLER_113_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14149_ net916 net695 VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__nand2_1
XFILLER_113_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18957_ _09840_ _09843_ _09845_ _09771_ VGND VGND VPWR VPWR _09849_ sky130_fd_sc_hd__o211ai_2
X_17908_ _08699_ _08735_ _08740_ VGND VGND VPWR VPWR _08767_ sky130_fd_sc_hd__o21ai_1
XFILLER_67_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18888_ net760 net596 net1001 net942 VGND VGND VPWR VPWR _09780_ sky130_fd_sc_hd__nand4_4
X_17839_ _08697_ _08699_ VGND VGND VPWR VPWR _08700_ sky130_fd_sc_hd__nand2_1
Xrebuffer25 net819 VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__buf_1
Xrebuffer14 b_l\[4\] VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer36 _00662_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__buf_6
Xrebuffer47 net843 VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer58 net648 VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer69 net861 VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_19_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20781_ clknet_leaf_19_clk _00421_ VGND VGND VPWR VPWR a_l\[3\] sky130_fd_sc_hd__dfxtp_4
X_19509_ _00692_ _00695_ _00588_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__o21ai_2
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer104 a_l\[11\] VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer137 net932 VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer115 a_h\[14\] VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__buf_8
XFILLER_135_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer159 a_h\[9\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer148 _06003_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd1_1
Xhold530 _00177_ VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap260 _06850_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_1
Xhold552 p_hl\[24\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _10115_ VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 mid_sum\[13\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ _01440_ net214 _01441_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__a21o_1
Xmax_cap271 net272 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
Xmax_cap282 _07035_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_1
Xhold574 term_high\[61\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20146_ _01234_ _01317_ _01309_ _01314_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__o22ai_1
XFILLER_131_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20077_ _01287_ _01290_ _01306_ _01308_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__o211ai_1
XFILLER_100_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11850_ _02766_ _02767_ _02780_ _02782_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__o211ai_1
X_11781_ _02524_ _02650_ _02655_ _02714_ _02716_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__o2111ai_2
XTAP_TAPCELL_ROW_103_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _01806_ _01807_ _01816_ _01817_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__or4_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10732_ p_hl\[16\] p_lh\[16\] _01760_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a21o_1
XFILLER_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13520_ _04424_ _04426_ _04428_ net954 VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_45_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ _01693_ _01697_ _01699_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__nand3_1
X_13451_ _04353_ _04357_ _04358_ _04344_ _04343_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__o2111ai_2
XFILLER_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16170_ _06952_ _07041_ _07042_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__nand3_2
X_10594_ net794 net1180 VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__and2_1
X_12402_ _03194_ _03197_ _03331_ _03332_ VGND VGND VPWR VPWR _03335_ sky130_fd_sc_hd__nand4_1
X_13382_ _04289_ _04285_ _04282_ _04290_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__o211ai_4
X_12333_ _09482_ _09613_ _03128_ _03261_ _03260_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__o221ai_4
X_15121_ net730 net657 VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__nand2_1
XFILLER_147_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15052_ _05946_ _05948_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__nand2_1
XFILLER_147_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ _03194_ _03195_ net398 VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__a21o_1
XFILLER_5_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14003_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__inv_2
X_11215_ net681 net525 net1052 net967 VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__a22oi_1
X_12195_ net906 net511 net508 net661 VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__a22oi_1
X_19860_ _00961_ _00964_ _00962_ VGND VGND VPWR VPWR _01077_ sky130_fd_sc_hd__a21o_1
Xoutput94 net94 VGND VGND VPWR VPWR p[35] sky130_fd_sc_hd__buf_2
X_11146_ _01857_ _02082_ _02078_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__o21ai_1
Xoutput72 net72 VGND VGND VPWR VPWR p[15] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18811_ net299 _09700_ net1031 net1081 VGND VGND VPWR VPWR _09704_ sky130_fd_sc_hd__o211ai_2
X_19791_ _00887_ _00882_ _00885_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__o21ai_4
Xoutput83 net83 VGND VGND VPWR VPWR p[25] sky130_fd_sc_hd__buf_2
X_15954_ _06825_ _06822_ _06742_ _06828_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__o211ai_4
X_11077_ net691 net1109 net1052 net697 VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__a22oi_1
X_18742_ _09626_ _09627_ _09628_ VGND VGND VPWR VPWR _09629_ sky130_fd_sc_hd__and3_1
XFILLER_49_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14905_ _05681_ _05797_ net745 net649 _05796_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__o2111ai_2
X_15885_ _06760_ _06762_ net1117 net541 VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__nand4_2
X_18673_ _09545_ _09549_ _09551_ _09547_ VGND VGND VPWR VPWR _09554_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_19_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17624_ _08486_ _08487_ VGND VGND VPWR VPWR _08488_ sky130_fd_sc_hd__nand2_2
XFILLER_64_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14836_ _05606_ _05607_ _05625_ _05621_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__a31o_1
X_17555_ _08413_ _08417_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__nand2_1
X_14767_ net716 net699 _05545_ _05543_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__a31o_1
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16506_ _07376_ _07378_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__nand2_1
X_11979_ _02891_ _02908_ _02744_ _02881_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__o2bb2ai_2
X_13718_ _04529_ _04540_ _04623_ _04622_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__o211ai_2
X_17486_ _08350_ _08351_ _08341_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__a21oi_2
X_14698_ _05475_ _05486_ _05487_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16437_ _07286_ _07221_ _07285_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__a21boi_2
XFILLER_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13649_ net714 net963 _04554_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__a31o_1
X_19225_ _09759_ _09902_ _09901_ VGND VGND VPWR VPWR _10123_ sky130_fd_sc_hd__o21ai_2
X_16368_ net1004 net1105 net523 net583 VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__a22oi_2
X_19156_ _10044_ _10045_ _10041_ VGND VGND VPWR VPWR _10048_ sky130_fd_sc_hd__a21oi_1
X_18107_ net458 _06401_ VGND VGND VPWR VPWR _08955_ sky130_fd_sc_hd__nand2_1
X_19087_ _09744_ net411 _09766_ _09768_ VGND VGND VPWR VPWR _09978_ sky130_fd_sc_hd__a22oi_2
X_15319_ _06212_ _06074_ _06213_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__a21oi_4
X_16299_ _06851_ _07043_ _07046_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__o21ai_2
X_18038_ _08886_ _08887_ net805 _06402_ VGND VGND VPWR VPWR _08888_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_141_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20000_ _01219_ _01223_ _09308_ _09319_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_140_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19989_ net731 net563 VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20764_ clknet_leaf_1_clk _00404_ VGND VGND VPWR VPWR a_h\[2\] sky130_fd_sc_hd__dfxtp_4
XFILLER_50_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20695_ clknet_leaf_4_clk _00335_ VGND VGND VPWR VPWR p_hl\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire718 b_l\[14\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__buf_6
XFILLER_6_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_131_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold360 p_hh\[0\] VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold371 p_ll_pipe\[4\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 p_hh\[3\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ net697 net519 VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__nand2_1
Xhold382 p_ll\[8\] VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
X_20129_ _01359_ _01363_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__nand2_1
XFILLER_133_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12951_ _03719_ _03723_ _03866_ _03861_ VGND VGND VPWR VPWR _03878_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_5_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_116_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11902_ net692 net489 VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__nand2_1
X_15670_ net309 _06533_ _06546_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__nand3_4
X_12882_ net659 b_h\[13\] VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__nand2_1
XFILLER_46_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11833_ net698 net487 VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nand2_1
X_14621_ _05521_ _05412_ _05522_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__nand3_2
X_17340_ net554 net514 VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__nand2_1
XFILLER_61_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11764_ _02524_ _02650_ _02655_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__o21a_1
X_14552_ _05452_ _05453_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__nand2_1
X_11695_ net664 net658 net526 net1059 _02626_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__a41o_1
X_17271_ _08133_ _08132_ _07993_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__nand3_4
X_10715_ p_hl\[13\] p_lh\[13\] _01748_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o21a_1
X_13503_ net789 net666 VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__nand2_1
X_14483_ _05223_ _05380_ _05381_ _05379_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__a31oi_1
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16222_ net572 net532 VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__nand2_1
X_10646_ net797 _01689_ _01690_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__nor3_1
X_13434_ _04343_ _04344_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__nand2_2
X_19010_ _09893_ _09897_ _09896_ _09871_ VGND VGND VPWR VPWR _09901_ sky130_fd_sc_hd__o211ai_4
XFILLER_42_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16153_ _09166_ _09646_ _07027_ _07028_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__o22a_2
Xrebuffer5 net801 VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd1_1
X_10577_ net795 net1274 VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_125_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13365_ _04274_ net705 net763 _04272_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_58_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15104_ net745 net640 net635 net750 VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__a22oi_2
X_12316_ _03112_ _03113_ _03123_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__a21oi_1
X_16084_ _06901_ _06958_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__nand2_2
XFILLER_127_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13296_ _04156_ _04176_ _04174_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__o21a_1
XFILLER_5_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ _03177_ _03179_ _03178_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_47_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19912_ _01126_ _01129_ _01125_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__a21oi_1
X_15035_ _05928_ _05930_ _05925_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a21oi_1
XFILLER_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19843_ _00939_ _00943_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__nand3_4
X_12178_ _02949_ _02952_ _02695_ _02955_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__a2bb2o_2
X_16986_ _07621_ _07853_ _07854_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__nand3_1
X_11129_ _02066_ _02068_ _02063_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__a21o_1
XFILLER_95_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19774_ net877 net820 net1102 net548 VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__nand4_2
XPHY_EDGE_ROW_134_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15937_ _06808_ _06809_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__nor2_1
X_18725_ net447 _09607_ _09609_ VGND VGND VPWR VPWR _09610_ sky130_fd_sc_hd__o21ai_1
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15868_ _09166_ _09624_ _06744_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__or3_1
XFILLER_64_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18656_ net618 net743 VGND VGND VPWR VPWR _09535_ sky130_fd_sc_hd__nand2_1
X_17607_ _08467_ _08469_ _08415_ VGND VGND VPWR VPWR _08471_ sky130_fd_sc_hd__nand3b_2
XTAP_TAPCELL_ROW_69_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14819_ net740 net736 net668 net663 VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__nand4_4
XFILLER_24_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15799_ net607 net527 VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__nand2_1
X_18587_ _09199_ _09264_ _09455_ _09456_ VGND VGND VPWR VPWR _09459_ sky130_fd_sc_hd__o211ai_2
X_17538_ _09297_ _09646_ _08397_ _08399_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_82_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17469_ _08179_ _08190_ _08328_ _08330_ VGND VGND VPWR VPWR _08335_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_43_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19208_ _10075_ _10100_ _10101_ VGND VGND VPWR VPWR _10105_ sky130_fd_sc_hd__and3_1
X_20480_ clknet_leaf_45_clk _00120_ VGND VGND VPWR VPWR term_mid\[24\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_143_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19139_ _10025_ _10020_ _10027_ _10010_ VGND VGND VPWR VPWR _10031_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_113_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20747_ clknet_leaf_42_clk _00387_ VGND VGND VPWR VPWR p_ll\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10500_ _01653_ net1331 term_high\[52\] VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__and3_1
Xwire515 net516 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_12
X_11480_ _02414_ _02415_ _02389_ _02390_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__o211ai_1
Xwire526 b_h\[3\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_8
X_20678_ clknet_leaf_55_clk _00318_ VGND VGND VPWR VPWR p_hl\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_7_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10431_ _01597_ _01598_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__nor2_1
Xwire559 a_l\[13\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__buf_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13150_ _03966_ _04009_ _04042_ _04044_ _04046_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__a221oi_1
X_10362_ term_low\[31\] term_mid\[31\] VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__nor2_1
XFILLER_136_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12101_ _02917_ _02969_ _03029_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__a21oi_1
XFILLER_88_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13081_ _03959_ _04002_ a_h\[12\] net478 _04004_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__o2111ai_2
X_10293_ term_low\[21\] term_mid\[21\] VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__nor2_1
X_12032_ _02937_ _02946_ _02936_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__a21boi_1
XFILLER_88_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_105_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16840_ _07707_ _07709_ net629 net472 VGND VGND VPWR VPWR _07711_ sky130_fd_sc_hd__and4_1
XFILLER_78_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16771_ net554 net1037 VGND VGND VPWR VPWR _07642_ sky130_fd_sc_hd__nand2_2
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13983_ _04744_ _04745_ _04743_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_144_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15722_ net607 net531 VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__nand2_1
X_12934_ _03775_ _03725_ _03774_ _03859_ _03860_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__o2111ai_2
X_18510_ _09155_ _09275_ net459 _07234_ _09374_ VGND VGND VPWR VPWR _09376_ sky130_fd_sc_hd__o221ai_4
XFILLER_46_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _00452_ _00477_ _00479_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__nand3_2
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15653_ net628 net515 VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__and2_1
X_12865_ _03791_ _03793_ _03790_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__o21ai_1
X_18441_ _09290_ _09295_ net252 _09296_ VGND VGND VPWR VPWR _09301_ sky130_fd_sc_hd__o211ai_2
XTAP_TAPCELL_ROW_29_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _06464_ _06465_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__nand2_1
X_11816_ _02721_ _02750_ _02751_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__nand3_4
X_12796_ _03718_ _03723_ _03722_ VGND VGND VPWR VPWR _03725_ sky130_fd_sc_hd__o21ai_2
X_18372_ _09223_ _09224_ VGND VGND VPWR VPWR _09225_ sky130_fd_sc_hd__nor2_1
X_14604_ _05414_ _05502_ _05503_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__nand3_2
XFILLER_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11747_ _02347_ _02467_ _02470_ _02677_ _02679_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__o2111ai_1
X_17323_ _08189_ VGND VGND VPWR VPWR _08190_ sky130_fd_sc_hd__inv_2
X_14535_ _05433_ net313 VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__nand2_1
X_17254_ net342 _08116_ _08101_ VGND VGND VPWR VPWR _08122_ sky130_fd_sc_hd__a21o_1
X_16205_ net973 net484 _07074_ _07076_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__a22o_1
X_11678_ _02608_ _02614_ VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__nand2_1
X_14466_ _05138_ _05356_ _05357_ _05220_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__a31o_1
X_10629_ p_hl\[1\] p_lh\[1\] VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__nand2_1
X_17185_ net558 net964 net969 net566 VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__a22oi_1
X_13417_ net435 _04324_ _04325_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__and3_1
X_14397_ _05147_ _05152_ _05150_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16136_ _06979_ _06987_ _06988_ _07006_ _07008_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__a32oi_4
X_13348_ net758 net753 VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__nand2_8
X_16067_ _06940_ _06943_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__nand2_1
X_13279_ net784 net693 net986 net787 VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__a22oi_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15018_ _05812_ _05813_ _05673_ _05914_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__a31o_2
XFILLER_142_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_130_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19826_ _00927_ _00937_ _01036_ _01037_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__a22oi_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19757_ _00725_ _00727_ _00961_ _00963_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__nand4_2
X_16969_ _07800_ _07801_ _07832_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__o21ai_2
X_18708_ _09588_ _09591_ net794 VGND VGND VPWR VPWR _09593_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19688_ _00882_ _00884_ _00886_ _00890_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__o31ai_1
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18639_ _09475_ _09516_ VGND VGND VPWR VPWR _09517_ sky130_fd_sc_hd__nand2_2
X_20601_ clknet_leaf_13_clk _00241_ VGND VGND VPWR VPWR p_hh_pipe\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20532_ clknet_leaf_47_clk _00172_ VGND VGND VPWR VPWR term_low\[27\] sky130_fd_sc_hd__dfxtp_1
X_20463_ clknet_leaf_14_clk _00103_ VGND VGND VPWR VPWR term_high\[55\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_118_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20394_ clknet_leaf_42_clk _00034_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10980_ _01920_ _01922_ _01917_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__a21o_1
XFILLER_83_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12650_ _03412_ _03413_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__nand2_1
XFILLER_70_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11601_ _02537_ _02539_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__nand2_2
X_12581_ _09504_ _09613_ _03509_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__o21ai_2
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14320_ _05218_ _05023_ _05217_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__nand3_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ _02467_ _02469_ _02347_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire312 _05563_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_4
XFILLER_139_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11463_ _02255_ net1018 net967 VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__nand3_1
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14251_ _05153_ _05154_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__nor2_2
X_10414_ _01574_ _01580_ _01581_ _01582_ _01584_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__o41a_2
Xwire378 _07648_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_1
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13202_ _04070_ _04085_ _04111_ _04109_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__o31a_1
Xwire367 _00752_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_1
X_14182_ _04864_ _04866_ _04862_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__a21o_1
X_11394_ _02334_ _02332_ net796 VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__a21o_1
XFILLER_125_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13133_ _04049_ _04055_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__nand3_1
X_18990_ _09749_ _09754_ _09752_ VGND VGND VPWR VPWR _09881_ sky130_fd_sc_hd__a21oi_1
X_10345_ _01106_ _01161_ net794 VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__o21ai_1
XFILLER_140_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_124_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17941_ _08786_ _08779_ _08785_ VGND VGND VPWR VPWR _08798_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13064_ _03957_ _03988_ _03989_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__nand3b_1
X_10276_ _10126_ _10137_ VGND VGND VPWR VPWR _10158_ sky130_fd_sc_hd__nor2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12015_ _02943_ _02944_ _02936_ _02937_ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__o211ai_1
X_17872_ _08730_ _08731_ _08724_ VGND VGND VPWR VPWR _08732_ sky130_fd_sc_hd__o21ai_1
X_16823_ _07680_ _07686_ _07685_ _07664_ net278 VGND VGND VPWR VPWR _07694_ sky130_fd_sc_hd__o2111ai_4
X_19611_ _00805_ _00807_ _00796_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__and3_1
Xclone235 net489 VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__clkbuf_16
XFILLER_65_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16754_ _07620_ _07621_ _07622_ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__and3_1
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19542_ _09220_ _09373_ _10170_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__or3_1
Xclone268 _00454_ _00465_ _00466_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__nand3_4
X_13966_ _04736_ _04737_ _04756_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__o21a_1
X_16685_ _07552_ _07553_ _07490_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__nand3_4
X_15705_ net346 net309 _06533_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__a21boi_2
XTAP_TAPCELL_ROW_66_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12917_ _03732_ _03839_ _03840_ VGND VGND VPWR VPWR _03845_ sky130_fd_sc_hd__nand3_1
X_13897_ _04668_ _04797_ _04798_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__and3_1
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19473_ _00648_ _00659_ _00660_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__nand3_4
X_15636_ _09210_ _09581_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__nor2_1
X_12848_ _03774_ _03776_ _03725_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__a21o_1
X_18424_ _09137_ _09139_ _09277_ _09278_ VGND VGND VPWR VPWR _09282_ sky130_fd_sc_hd__o211ai_4
XTAP_TAPCELL_ROW_66_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ _06435_ _06447_ _06449_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__and3_1
X_12779_ _03697_ _03612_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__nand2_1
X_18355_ _09203_ _09200_ _09099_ _09201_ VGND VGND VPWR VPWR _09207_ sky130_fd_sc_hd__a211oi_4
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18286_ _09058_ _09074_ _09073_ _09071_ VGND VGND VPWR VPWR _09132_ sky130_fd_sc_hd__o2bb2ai_1
X_17306_ net573 net569 net498 net493 _08168_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__a41o_1
X_14518_ net756 net655 VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__nand2_1
X_15498_ net716 net635 _06369_ _06371_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17237_ net582 net493 VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__nand2_1
X_14449_ _09308_ _09428_ _05204_ _05347_ _05346_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__o221ai_4
XFILLER_30_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap601 net602 VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__buf_12
Xmax_cap612 a_l\[4\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__buf_8
X_17168_ _07967_ _07969_ _07978_ _07985_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__o211ai_2
X_16119_ net966 net515 VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__nand2_1
Xmax_cap623 net625 VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__buf_12
Xmax_cap645 a_h\[13\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_12
Xmax_cap634 a_h\[15\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__buf_12
XFILLER_6_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap678 net679 VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__buf_12
X_17099_ net608 net600 net485 net479 VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__and4_1
Xmax_cap656 net657 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__buf_8
Xmax_cap667 net669 VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__buf_12
XFILLER_142_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_115_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap689 net690 VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__buf_8
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19809_ _01017_ _01018_ _01020_ _00915_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_28_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20515_ clknet_leaf_41_clk _00155_ VGND VGND VPWR VPWR term_low\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_20446_ clknet_leaf_27_clk _00086_ VGND VGND VPWR VPWR term_high\[38\] sky130_fd_sc_hd__dfxtp_1
XFILLER_118_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20377_ clknet_leaf_35_clk _00017_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfxtp_1
XFILLER_133_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_141_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13820_ _04718_ _04725_ _04724_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__o21ai_2
XFILLER_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10963_ net702 net1052 VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__nand2_1
XFILLER_62_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13751_ _04586_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__nand2_1
XFILLER_44_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16470_ _07338_ _07341_ _07340_ VGND VGND VPWR VPWR _07343_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_106_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12702_ _03628_ _03629_ _09449_ _09668_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_48_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13682_ _04518_ _04520_ _04522_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__o21ai_1
X_10894_ net794 net1160 VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__and2_1
X_15421_ _06310_ _06311_ _09362_ _09515_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__o2bb2a_1
X_12633_ _03535_ _03558_ _03560_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__nor3_1
XTAP_TAPCELL_ROW_139_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _03492_ _03494_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__nand2_1
X_18140_ _08984_ _08985_ VGND VGND VPWR VPWR _08988_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_61_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ _06000_ _06178_ _06242_ _06186_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__o211ai_2
XFILLER_8_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11515_ net698 net497 VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__nand2_1
X_18071_ _08917_ _08918_ VGND VGND VPWR VPWR _08920_ sky130_fd_sc_hd__nand2_2
X_15283_ _06172_ _06176_ _06177_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__o21ai_1
X_14303_ net736 net685 VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__nand2_2
XFILLER_144_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17022_ _07888_ _07889_ _07770_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__and3b_1
X_12495_ _03278_ _03281_ _03280_ VGND VGND VPWR VPWR _03427_ sky130_fd_sc_hd__o21ai_2
X_14234_ _05120_ _05134_ _05136_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__a21boi_2
XFILLER_109_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11446_ _02370_ _02372_ _02379_ _02381_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__nand4_1
Xwire197 _04316_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11377_ _02246_ _02247_ _02315_ _02316_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__a22o_1
X_14165_ _05050_ _05066_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__nand2_1
X_13116_ _04033_ _04038_ _04040_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__a21oi_1
X_18973_ _09863_ _09864_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__nor2_1
X_14096_ _04994_ _04997_ net392 VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a21o_1
X_10328_ _00870_ _00978_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__nand2_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17924_ _09373_ _09668_ _08781_ VGND VGND VPWR VPWR _08782_ sky130_fd_sc_hd__or3_1
X_13047_ _03962_ _03963_ _03970_ _03971_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__nand4_2
X_10259_ net794 net1250 VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__and2_1
X_17855_ _08715_ _08712_ VGND VGND VPWR VPWR _08716_ sky130_fd_sc_hd__nand2_1
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16806_ _07670_ _07672_ _07667_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__a21o_1
X_17786_ _09297_ _09657_ _08553_ _08558_ VGND VGND VPWR VPWR _08648_ sky130_fd_sc_hd__o31a_1
X_16737_ _07604_ _07605_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__nand2_1
X_19525_ net797 _00715_ _00716_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__nor3b_1
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14998_ _05835_ _05836_ _05839_ _05850_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__o2111ai_4
XFILLER_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13949_ _04850_ _04853_ _04849_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__o21ai_1
X_16668_ _07520_ _07539_ VGND VGND VPWR VPWR _07540_ sky130_fd_sc_hd__nand2_2
XFILLER_61_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19456_ _00640_ _00641_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__nor2_1
X_16599_ net620 net484 net480 net840 VGND VGND VPWR VPWR _07471_ sky130_fd_sc_hd__a22oi_2
X_15619_ _06455_ _06459_ _06499_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__nand3_1
X_18407_ _09257_ _09258_ _09243_ _09247_ VGND VGND VPWR VPWR _09263_ sky130_fd_sc_hd__o211ai_2
XFILLER_61_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19387_ _00561_ _00562_ _00564_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18338_ net457 _06402_ net336 _09038_ VGND VGND VPWR VPWR _09189_ sky130_fd_sc_hd__o31a_1
XFILLER_147_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer319 net587 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_79_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18269_ net626 net749 VGND VGND VPWR VPWR _09115_ sky130_fd_sc_hd__nand2_1
X_20300_ _01532_ _01536_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__o21ba_1
Xmax_cap420 _07204_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_1
Xmax_cap453 _07391_ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__buf_4
XFILLER_115_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap442 _01779_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__buf_1
Xmax_cap431 _04792_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__buf_1
X_20231_ net1013 b_l\[15\] _01472_ _01473_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__a22o_1
Xmax_cap464 _02105_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_92_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap486 b_h\[12\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_8
Xmax_cap475 b_h\[14\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_6
X_20162_ _01338_ _01342_ _01399_ _01400_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a22o_1
Xmax_cap497 net499 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_12
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20093_ _01326_ _01327_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__nand2_1
XFILLER_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ _02219_ _02225_ _02216_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__a21boi_1
XFILLER_119_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12280_ _03172_ _03212_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__nand2_1
X_20429_ clknet_leaf_15_clk _00069_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11231_ _02169_ _02171_ _02165_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__a21o_1
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11162_ net702 net510 net507 net707 VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__a22oi_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15970_ _09624_ _09635_ _06402_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__or3_4
X_11093_ net983 net507 VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__nand2_1
XFILLER_76_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14921_ _05814_ _05815_ _05817_ _05701_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__o211ai_4
X_17640_ _08396_ _08402_ _08500_ VGND VGND VPWR VPWR _08504_ sky130_fd_sc_hd__o21ai_1
X_14852_ _05749_ _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__nand2_1
X_13803_ net757 net752 net689 net683 VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__nand4_1
X_11995_ _02925_ _02928_ _02858_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a21o_1
X_17571_ _08329_ _08434_ _08435_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__nand3_2
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_55_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14783_ _05681_ _05682_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__nand2_2
X_19310_ net298 _00452_ _00473_ _00475_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__nand4_4
X_10946_ _01891_ net1106 net702 _01889_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__nand4_2
X_16522_ _06878_ _07392_ _07390_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__o21ai_4
X_13734_ _04639_ _04640_ _04629_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__nand3_2
XFILLER_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16453_ net812 net928 net496 net491 VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__nand4_1
X_10877_ _09690_ net1185 VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__and2_1
X_13665_ _04391_ _04392_ _04572_ _04570_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__o22ai_4
X_19241_ _10136_ _10006_ _10135_ VGND VGND VPWR VPWR _10141_ sky130_fd_sc_hd__nand3_4
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16384_ _06961_ _07129_ _07133_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__o21ai_2
X_12616_ _03542_ _03543_ net436 VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__a21oi_1
X_15404_ _06295_ _06294_ _06291_ _06296_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__o2bb2ai_1
X_19172_ _10032_ _10060_ VGND VGND VPWR VPWR _10066_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18123_ net790 net781 net601 net594 VGND VGND VPWR VPWR _08971_ sky130_fd_sc_hd__nand4_2
X_13596_ _04428_ net954 _04427_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__a21boi_4
X_15335_ net730 net635 VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__nand2_1
XFILLER_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12547_ _03463_ _03464_ _03472_ _03474_ VGND VGND VPWR VPWR _03479_ sky130_fd_sc_hd__o2bb2ai_2
XANTENNA_3 _00054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_18054_ _08865_ _08880_ _08879_ VGND VGND VPWR VPWR _08903_ sky130_fd_sc_hd__o21ai_2
X_12478_ _03394_ _03395_ _03405_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__nand3_1
X_15266_ net730 net643 VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__nand2_1
XFILLER_8_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17005_ _07868_ _07869_ _07870_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__a21o_1
X_11429_ _02366_ _02368_ _02355_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__a21oi_2
X_14217_ _04973_ _04976_ _04974_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__a21oi_1
X_15197_ net733 net910 net641 net739 VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__a22oi_1
X_14148_ net740 net690 VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__nand2_2
XFILLER_113_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18956_ _09844_ _09845_ _09771_ VGND VGND VPWR VPWR _09848_ sky130_fd_sc_hd__a21o_1
X_14079_ net783 net643 VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__nand2_1
X_17907_ _08764_ _08727_ _08765_ VGND VGND VPWR VPWR _08766_ sky130_fd_sc_hd__a21o_1
X_18887_ _09777_ _09778_ VGND VGND VPWR VPWR _09779_ sky130_fd_sc_hd__nand2_1
XFILLER_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17838_ _08698_ _08694_ VGND VGND VPWR VPWR _08699_ sky130_fd_sc_hd__nand2_1
XFILLER_67_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer15 a_l\[4\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer26 b_h\[10\] VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 net843 VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd1_1
X_17769_ net1054 net484 net480 net566 VGND VGND VPWR VPWR _08631_ sky130_fd_sc_hd__a22o_1
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer59 b_h\[9\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer37 b_l\[9\] VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd1_1
Xclkbuf_leaf_46_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_8
X_20780_ clknet_leaf_20_clk _00420_ VGND VGND VPWR VPWR a_l\[2\] sky130_fd_sc_hd__dfxtp_4
X_19508_ _00586_ _00587_ _00685_ _00694_ _00693_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__o221ai_2
X_19439_ _00607_ _00608_ _00623_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer105 _03953_ VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer138 net932 VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer116 net912 VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_136_727 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer149 net945 VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold520 _00032_ VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold531 p_hh\[28\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap250 _01483_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
X_20214_ _01451_ _01455_ _01456_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__a21oi_1
Xhold542 mid_sum\[14\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 term_mid\[23\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold575 term_high\[59\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap294 _02994_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold564 p_lh\[29\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_106_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20145_ _01312_ _01313_ _01101_ _01318_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__a31o_1
XFILLER_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_20076_ _01306_ _01308_ _01292_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__a21oi_2
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_37_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_8
X_11780_ _02651_ _02655_ _02714_ _02716_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ p_hl\[25\] p_lh\[25\] _01806_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__a21oi_1
X_10731_ p_hl\[17\] p_lh\[17\] VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_45_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13450_ _04343_ _04344_ _04359_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nand3_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ _03194_ _03197_ _03331_ _03332_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__a22o_1
X_10662_ p_hl\[6\] p_lh\[6\] VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__nor2_1
XFILLER_9_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10593_ net793 net1319 VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__and2_1
X_13381_ _04289_ _04285_ _04282_ _04290_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__o211a_1
X_12332_ _03128_ _03261_ net1019 b_h\[8\] _03260_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__o2111ai_4
X_15120_ _05925_ _05929_ _05928_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__o21a_1
X_12263_ net398 _03195_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nand2_2
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15051_ _05945_ _05947_ VGND VGND VPWR VPWR _05949_ sky130_fd_sc_hd__nor2_1
XFILLER_31_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11214_ net681 net525 VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__nand2_1
X_14002_ _04884_ _04885_ _04904_ _04906_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__o211ai_4
XFILLER_134_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12194_ net653 net511 VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__nand2_2
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11145_ _01857_ _02082_ _02078_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__o21a_1
XFILLER_96_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput73 net73 VGND VGND VPWR VPWR p[16] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18810_ _09697_ _09700_ _09676_ VGND VGND VPWR VPWR _09703_ sky130_fd_sc_hd__o21ai_1
Xoutput84 net84 VGND VGND VPWR VPWR p[26] sky130_fd_sc_hd__buf_2
XFILLER_1_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19790_ _00885_ _00887_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__nand2_1
Xoutput95 net95 VGND VGND VPWR VPWR p[36] sky130_fd_sc_hd__buf_2
X_15953_ _06742_ _06828_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__nand2_1
X_11076_ net691 net525 VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__nand2_1
X_18741_ net630 net729 _09544_ _09545_ VGND VGND VPWR VPWR _09628_ sky130_fd_sc_hd__a31o_1
XFILLER_1_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14904_ _05681_ _05797_ _05800_ _05796_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__o211a_4
X_15884_ net602 net595 net531 net527 VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__nand4_4
X_18672_ _09547_ _09550_ _09551_ VGND VGND VPWR VPWR _09553_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_91_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17623_ net581 net476 _08483_ _08484_ VGND VGND VPWR VPWR _08487_ sky130_fd_sc_hd__a22o_1
XFILLER_63_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14835_ _05565_ _05580_ _05583_ _05729_ _05730_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__o2111ai_1
X_11978_ net323 _02907_ _02891_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__a21o_1
XFILLER_91_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17554_ _08416_ _08418_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__nand2_1
X_14766_ _09690_ _05665_ _05666_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__and3_1
X_10929_ _01875_ _01876_ _01866_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__a21oi_1
X_16505_ net570 net561 net533 net529 VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__nand4_4
XFILLER_72_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13717_ _04621_ _04588_ _04620_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nand3_4
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17485_ _08231_ _08234_ _08339_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__o21ai_2
X_19224_ net1128 net718 _09873_ _09874_ VGND VGND VPWR VPWR _10122_ sky130_fd_sc_hd__a31o_1
X_14697_ _05589_ _05458_ _05590_ _05594_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__nand4_4
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16436_ _07285_ _07287_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__nand2_1
X_13648_ net714 net734 net963 net741 VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__a22oi_2
XFILLER_32_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16367_ _07236_ _07237_ _07227_ VGND VGND VPWR VPWR _07241_ sky130_fd_sc_hd__nand3_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13579_ _01871_ _04260_ _04446_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__o21ai_2
XFILLER_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19155_ _10045_ _10044_ net765 net568 VGND VGND VPWR VPWR _10047_ sky130_fd_sc_hd__and4_1
X_16298_ _06951_ _07038_ _07040_ _06851_ VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__a31oi_2
XFILLER_118_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18106_ _08933_ _08931_ _08900_ _08938_ VGND VGND VPWR VPWR _08954_ sky130_fd_sc_hd__a22oi_2
X_19086_ _09869_ _09972_ _09973_ VGND VGND VPWR VPWR _09977_ sky130_fd_sc_hd__nand3_4
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15318_ _06079_ _06140_ _06141_ _06071_ _06144_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__a32o_1
X_18037_ _08857_ _08882_ _08883_ VGND VGND VPWR VPWR _08887_ sky130_fd_sc_hd__nand3b_2
X_15249_ _06140_ _06141_ _06079_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__nand3_1
XFILLER_125_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19988_ _01211_ _01208_ _01213_ VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__a21oi_4
XFILLER_101_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18939_ _09807_ _09824_ VGND VGND VPWR VPWR _09831_ sky130_fd_sc_hd__nand2_1
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20763_ clknet_leaf_1_clk _00403_ VGND VGND VPWR VPWR a_h\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20694_ clknet_leaf_4_clk _00334_ VGND VGND VPWR VPWR p_hl\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire719 net720 VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__buf_6
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold361 p_hh\[4\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold394 p_hh_pipe\[31\] VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 p_ll_pipe\[0\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 p_ll\[23\] VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
X_20128_ _01218_ _01361_ _01362_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__o21ai_1
XFILLER_131_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_133_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12950_ _03875_ _03876_ _03877_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_5_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ net574 net721 _01285_ _01286_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__a22o_1
X_11901_ net687 net682 net497 net492 VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__nand4_4
XFILLER_93_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12881_ net396 _03756_ _03754_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__a21boi_2
XFILLER_46_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11832_ _01888_ _02338_ _02578_ _02579_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__o22ai_4
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14620_ _05508_ _05518_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__nand2_1
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14551_ _04987_ _05285_ _05448_ _05449_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__o211ai_2
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11763_ _02664_ _02644_ _02642_ _02645_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__o2bb2ai_1
X_11694_ net462 _02629_ _02626_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__o21ai_2
X_17270_ _08083_ _08136_ _08134_ _07992_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__o211ai_4
X_10714_ _01736_ _01740_ _01743_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__nand3b_2
X_13502_ net785 net673 VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__nand2_1
X_14482_ _01871_ net455 _05195_ _05224_ _05382_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__o2111ai_4
X_16221_ net582 net528 VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__nand2_1
X_10645_ _01680_ _01684_ _01688_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__a21boi_1
X_13433_ _04338_ _04342_ _04336_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16152_ net841 net629 net496 net491 VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__and4_1
X_13364_ _04272_ net705 net763 VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__and3_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_850 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12315_ _03244_ _03248_ _03247_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__o21ai_1
XFILLER_127_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer6 net800 VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_58_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15103_ net751 net745 net914 net635 VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__nand4_4
X_10576_ _09690_ net1340 VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__and2_1
X_16083_ net607 net512 net505 net613 VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__a22oi_1
X_13295_ _04207_ _04204_ _04206_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__a21o_1
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12246_ _03177_ _03179_ _03178_ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__a21oi_1
XFILLER_5_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_19911_ _09275_ _09286_ _05044_ _01125_ _01126_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__o311a_1
X_15034_ _05930_ net663 net730 _05928_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__nand4_1
X_12177_ _03110_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_71_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19842_ _09231_ _09362_ _00904_ _00903_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__o31a_1
XFILLER_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11128_ _09406_ _09602_ _02020_ _02067_ _02066_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__o221ai_2
XFILLER_69_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16985_ _07621_ _07853_ _07854_ VGND VGND VPWR VPWR _07855_ sky130_fd_sc_hd__and3_1
XFILLER_95_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19773_ _00872_ _00982_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__nand2_1
X_15936_ _06789_ _06799_ _06800_ _06804_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__and4_1
X_11059_ net967 net534 VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__nand2_1
XFILLER_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18724_ net621 net732 VGND VGND VPWR VPWR _09609_ sky130_fd_sc_hd__nand2_2
X_15867_ _06743_ _06744_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__nor2_2
X_18655_ net621 net737 VGND VGND VPWR VPWR _09534_ sky130_fd_sc_hd__nand2_1
X_17606_ _08413_ _08467_ _08468_ VGND VGND VPWR VPWR _08470_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_69_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14818_ _05616_ _05716_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__nand2_1
X_15798_ net595 net541 VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__nand2_1
X_18586_ _09455_ _09456_ net610 net749 VGND VGND VPWR VPWR _09458_ sky130_fd_sc_hd__nand4_1
X_17537_ _09297_ _09646_ _08309_ _08395_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__o22a_1
X_14749_ _05546_ _05548_ _05641_ _05551_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__a22o_1
XFILLER_32_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17468_ _08329_ _08331_ _08301_ VGND VGND VPWR VPWR _08334_ sky130_fd_sc_hd__nand3_2
XTAP_TAPCELL_ROW_43_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16419_ _07289_ _07292_ VGND VGND VPWR VPWR _07293_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19207_ _10076_ _10102_ _10103_ VGND VGND VPWR VPWR _10104_ sky130_fd_sc_hd__nand3_1
XFILLER_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17399_ _08036_ _08038_ VGND VGND VPWR VPWR _08266_ sky130_fd_sc_hd__nand2_1
X_19138_ _10028_ _10009_ VGND VGND VPWR VPWR _10030_ sky130_fd_sc_hd__nand2_1
XFILLER_146_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_8_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_19069_ _09958_ _09959_ VGND VGND VPWR VPWR _09960_ sky130_fd_sc_hd__nand2_1
XFILLER_133_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_20746_ clknet_leaf_42_clk _00386_ VGND VGND VPWR VPWR p_ll\[16\] sky130_fd_sc_hd__dfxtp_1
X_10430_ term_mid\[41\] term_high\[41\] VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__and2_1
Xwire516 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_12
Xwire549 net550 VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__buf_8
X_20677_ clknet_leaf_55_clk _00317_ VGND VGND VPWR VPWR p_hl\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10361_ net471 _01322_ _01333_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__a21oi_1
XFILLER_124_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12100_ net1047 _02970_ _03031_ _03029_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__o2bb2ai_4
X_13080_ _09515_ _09657_ _04002_ _04004_ _04001_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__o311a_1
X_10292_ _00558_ _00579_ _00590_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__o21a_1
X_12031_ _02964_ _02965_ _02966_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__o21a_1
XFILLER_105_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16770_ net558 net530 VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__nand2_1
X_13982_ _04876_ _04883_ _04886_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_144_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ net1090 net527 VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__nand2_1
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12933_ _03775_ _03725_ _03774_ _03859_ _03860_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__o2111a_1
X_18440_ _09298_ _09225_ VGND VGND VPWR VPWR _09300_ sky130_fd_sc_hd__nand2_1
XFILLER_46_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15652_ _06523_ _06529_ _06515_ _06531_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__o211ai_4
X_12864_ _03605_ net136 _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ net607 net542 VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__nand2_1
X_11815_ _02749_ _02720_ _02748_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__nand3_4
X_12795_ _03719_ _03720_ _03716_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__and3_1
X_18371_ _09124_ _09128_ _09219_ VGND VGND VPWR VPWR _09224_ sky130_fd_sc_hd__and3_1
XFILLER_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14603_ _05465_ _05499_ _05501_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__nand3_1
X_11746_ _02677_ _02679_ _02681_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__a21bo_1
X_17322_ _08177_ net341 _08184_ _08186_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__nand4_4
X_14534_ _05305_ _05431_ _05430_ _05428_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__o211a_1
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17253_ net342 _08116_ _08101_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__nand3_2
X_16204_ _07074_ _07076_ net973 net484 VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__nand4_1
XFILLER_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11677_ _02612_ _02614_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_40_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14465_ _05138_ _05356_ _05357_ _05220_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__a31oi_2
X_10628_ p_hl\[1\] p_lh\[1\] VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__and2_1
X_17184_ net559 net514 VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__nand2_4
X_13416_ net435 _04324_ _04325_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__a21o_1
X_14396_ _05147_ _05152_ _05150_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__a21o_1
X_10559_ net793 net1288 VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__and2_1
X_16135_ _06990_ _06994_ _07002_ _07003_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__o2bb2ai_2
X_13347_ net753 net758 VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__and2_4
X_16066_ _06826_ _06831_ _06729_ _06834_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__o22ai_1
X_13278_ net777 net700 VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__nand2_1
X_12229_ net357 _03023_ _03157_ _03159_ VGND VGND VPWR VPWR _03163_ sky130_fd_sc_hd__nand4_4
X_15017_ _05911_ _05912_ _05811_ _05816_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__o22a_1
XFILLER_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_19825_ _00927_ _00937_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__nand2_1
XFILLER_111_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16968_ _07805_ _07830_ _07831_ VGND VGND VPWR VPWR _07838_ sky130_fd_sc_hd__nand3_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_19756_ _00725_ _00727_ _00961_ _00963_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__a22o_1
X_15919_ net617 net505 VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__nand2_1
X_18707_ _09313_ _09436_ _09440_ _09322_ VGND VGND VPWR VPWR _09591_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_37_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16899_ _07743_ _07745_ _07760_ _07762_ VGND VGND VPWR VPWR _07769_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_84_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19687_ _00881_ _00886_ net407 VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__a21oi_1
X_18638_ net301 _09496_ _09503_ net370 VGND VGND VPWR VPWR _09516_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_37_577 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18569_ _09313_ _09436_ _09440_ VGND VGND VPWR VPWR _09441_ sky130_fd_sc_hd__a21o_1
X_20600_ clknet_leaf_12_clk _00240_ VGND VGND VPWR VPWR p_hh_pipe\[30\] sky130_fd_sc_hd__dfxtp_1
X_20531_ clknet_leaf_47_clk _00171_ VGND VGND VPWR VPWR term_low\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20462_ clknet_leaf_14_clk _00102_ VGND VGND VPWR VPWR term_high\[54\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_115_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20393_ clknet_leaf_37_clk _00033_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfxtp_1
XFILLER_134_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_114_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11600_ _02399_ _02402_ _02532_ _02533_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__nand4_1
X_12580_ _03506_ _03508_ net647 b_h\[8\] VGND VGND VPWR VPWR _03511_ sky130_fd_sc_hd__nand4_2
X_11531_ _02464_ _02466_ _02465_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__nand3_1
XFILLER_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20729_ clknet_leaf_6_clk _00369_ VGND VGND VPWR VPWR p_lh\[31\] sky130_fd_sc_hd__dfxtp_1
Xwire302 _09469_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__buf_1
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11462_ _02256_ _02397_ _02393_ _02396_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__o211ai_2
XFILLER_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14250_ _02502_ _04182_ net761 net662 _05151_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__o2111a_4
X_10413_ net796 _01583_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__nor2_1
X_11393_ _02143_ _02236_ _02147_ _02333_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__o22ai_4
X_13201_ _04107_ _04108_ _04070_ _04085_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__o2bb2a_1
X_14181_ _05082_ net210 net195 VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__a21o_1
Xwire368 _09912_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_1
XFILLER_125_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13132_ _09504_ _09679_ _04053_ _04054_ VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__o211ai_1
X_10344_ _00988_ _01150_ _01128_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__a21oi_2
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17940_ net555 a_l\[15\] net477 net473 _08796_ VGND VGND VPWR VPWR _08797_ sky130_fd_sc_hd__a41o_1
X_13063_ _03931_ _03932_ _03986_ _03987_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__nand4_1
X_10275_ term_low\[18\] term_mid\[18\] VGND VGND VPWR VPWR _10148_ sky130_fd_sc_hd__nand2_1
X_12014_ _02936_ _02937_ _02946_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__a21o_1
X_17871_ _08726_ _08727_ a_l\[12\] net473 VGND VGND VPWR VPWR _08731_ sky130_fd_sc_hd__and4_1
XFILLER_120_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16822_ _07664_ net278 _07684_ _07687_ VGND VGND VPWR VPWR _07693_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_19610_ _00808_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__inv_2
XFILLER_93_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19541_ net919 net765 net552 net548 VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__and4_2
X_16753_ _07620_ _07621_ _07622_ VGND VGND VPWR VPWR _07624_ sky130_fd_sc_hd__a21oi_1
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13965_ _04727_ _04767_ _04762_ _04764_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__o2bb2ai_1
X_16684_ _07552_ _07553_ _07490_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__and3_1
X_15704_ net387 _06583_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__nor2_8
X_12916_ _03842_ net397 _03841_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__nand3_2
X_13896_ _04797_ _04798_ _04667_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__a21o_1
X_19472_ _00654_ _00656_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__nand2_1
X_15635_ _06479_ _06486_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__nand2_1
X_12847_ _03772_ _03773_ _03727_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a21o_1
X_18423_ _09137_ _09139_ _09277_ _09278_ VGND VGND VPWR VPWR _09281_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _09202_ _09204_ _09099_ VGND VGND VPWR VPWR _09206_ sky130_fd_sc_hd__a21boi_1
X_12778_ _03704_ _03706_ _03707_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__a21oi_1
X_15566_ _06443_ _06445_ net423 VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__o21bai_2
X_17305_ net449 _08170_ _08168_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__o21ai_1
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11729_ _02644_ _02647_ _02664_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__nand3_2
X_18285_ _09129_ _09130_ VGND VGND VPWR VPWR _09131_ sky130_fd_sc_hd__nand2_1
X_15497_ _06385_ _06364_ net795 _06386_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__o211a_1
X_14517_ net750 net662 VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nand2_1
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17236_ net585 net488 VGND VGND VPWR VPWR _08104_ sky130_fd_sc_hd__nand2_1
X_14448_ _05346_ _05348_ _05343_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__a21o_1
Xmax_cap602 a_l\[6\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__buf_12
X_17167_ _07980_ _07981_ _08033_ _08034_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__o211ai_1
Xmax_cap624 net625 VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__buf_6
XFILLER_127_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap613 a_l\[4\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__buf_6
XFILLER_116_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16118_ _06992_ _06978_ _06991_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__nand3_2
X_14379_ _05280_ _05281_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__nand2_1
Xmax_cap635 net636 VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_8
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17098_ net600 net485 net479 net608 VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__a22oi_4
Xmax_cap679 net680 VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__buf_12
Xmax_cap646 net647 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_12
Xmax_cap657 a_h\[11\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkbuf_8
Xmax_cap668 net956 VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__clkbuf_8
X_16049_ _06921_ _06854_ _06919_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__nand3_2
XFILLER_131_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19808_ net742 net735 net567 net563 VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__nand4_1
XFILLER_84_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_19739_ _00810_ _00941_ _00940_ _00939_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__o211ai_2
XFILLER_38_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_20514_ clknet_leaf_31_clk _00154_ VGND VGND VPWR VPWR term_low\[9\] sky130_fd_sc_hd__dfxtp_1
X_20445_ clknet_leaf_27_clk _00085_ VGND VGND VPWR VPWR term_high\[37\] sky130_fd_sc_hd__dfxtp_1
XFILLER_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_106_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_20376_ clknet_leaf_35_clk _00016_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ net702 net1109 net519 net707 VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__a22oi_2
XFILLER_90_428 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13750_ _04625_ net287 _04643_ _04645_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12701_ _03629_ net475 net680 _03628_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__nand4_2
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13681_ net777 net673 _04416_ _04519_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__o2bb2a_2
X_10893_ net794 net1192 VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__and2_1
X_15420_ _06310_ _06311_ net719 net643 VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__and4_1
X_12632_ _03558_ _03560_ _03535_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__o21ai_4
X_12563_ _03493_ _03489_ _03491_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a21oi_2
X_15351_ _06000_ _06178_ _06242_ _06186_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__o211a_1
XFILLER_8_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11514_ net706 net492 VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__nand2_1
Xwire132 net133 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__buf_1
X_18070_ net781 net605 net601 net790 VGND VGND VPWR VPWR _08919_ sky130_fd_sc_hd__a22oi_1
X_12494_ _03151_ _03279_ _03278_ VGND VGND VPWR VPWR _03426_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_61_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15282_ _06154_ _06156_ _06173_ _06175_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__a22o_1
XFILLER_8_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14302_ _05056_ _05204_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__nand2_2
X_17021_ _07740_ net377 _07770_ _07889_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__a22oi_4
X_11445_ _02370_ _02372_ _02378_ _02380_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire143 _01271_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
X_14233_ _05120_ _05134_ _05135_ _05132_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_109_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire176 _03478_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
Xwire187 _09093_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
XFILLER_137_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11376_ _02246_ _02247_ _02315_ _02316_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__nand4_1
XFILLER_124_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14164_ _05048_ _05049_ net350 _05066_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__nand4_1
XFILLER_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13115_ _04033_ _04038_ net793 VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__o21ai_1
X_18972_ _09730_ _09735_ _09862_ net797 VGND VGND VPWR VPWR _09864_ sky130_fd_sc_hd__a31o_1
X_14095_ _04974_ _04977_ _04978_ _04998_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o211a_1
X_10327_ term_low\[24\] term_mid\[24\] _00902_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__a21oi_1
X_17923_ net473 _08676_ _08780_ net480 VGND VGND VPWR VPWR _08781_ sky130_fd_sc_hd__o22a_1
X_10258_ net794 net1194 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__and2_1
X_13046_ net394 _03963_ _03970_ _03971_ VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__a22o_1
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17854_ _08713_ _08624_ _08714_ VGND VGND VPWR VPWR _08715_ sky130_fd_sc_hd__o21bai_4
X_10189_ net592 VGND VGND VPWR VPWR _09242_ sky130_fd_sc_hd__inv_12
X_16805_ _09253_ _09613_ _07495_ _07671_ _07670_ VGND VGND VPWR VPWR _07676_ sky130_fd_sc_hd__o221ai_4
XFILLER_93_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17785_ a_l\[10\] net472 VGND VGND VPWR VPWR _08647_ sky130_fd_sc_hd__nand2_1
X_14997_ _05853_ _05856_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__nand2_1
X_16736_ net594 net498 net493 net600 VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__a22oi_2
X_19524_ _00707_ _00708_ _00714_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__nand3_1
XFILLER_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13948_ _04847_ _04848_ _04840_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__a21o_1
X_19455_ _00638_ _00639_ _00636_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__a21oi_2
XFILLER_35_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16667_ net379 _07536_ _07538_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__o21ai_1
X_18406_ _09243_ _09247_ _09252_ _09255_ VGND VGND VPWR VPWR _09262_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_62_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13879_ net731 net709 _04783_ _04784_ VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a22o_1
X_16598_ _07468_ _07469_ VGND VGND VPWR VPWR _07470_ sky130_fd_sc_hd__nand2_1
X_15618_ _06455_ _06459_ _06499_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__a21o_1
X_19386_ net216 _10121_ _10125_ _00561_ _00562_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__o2111ai_1
XTAP_TAPCELL_ROW_17_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15549_ net631 net522 VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__nand2_1
X_18337_ net630 net1082 VGND VGND VPWR VPWR _09187_ sky130_fd_sc_hd__nand2_2
X_18268_ _09048_ _09052_ _09049_ VGND VGND VPWR VPWR _09114_ sky130_fd_sc_hd__a21oi_4
XFILLER_147_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17219_ _07958_ _07960_ _07950_ _07974_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_79_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18199_ _08972_ _08981_ _08980_ _08994_ VGND VGND VPWR VPWR _09046_ sky130_fd_sc_hd__a2bb2oi_2
Xmax_cap443 _01590_ VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_1
Xmax_cap421 net422 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_1
X_20230_ _01472_ _01473_ _01469_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__a21oi_1
Xmax_cap454 _05160_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_4
XFILLER_143_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap487 net489 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_12
Xmax_cap465 _02080_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_92_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap476 net478 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_6
X_20161_ _01338_ _01342_ _01399_ _01400_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__a22oi_1
X_20092_ _01204_ _01207_ _01210_ _01244_ _01248_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__o2111ai_4
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_20428_ clknet_leaf_15_clk _00068_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_134_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ _09449_ _09592_ _02079_ _02170_ _02169_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__o221ai_4
XFILLER_106_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11161_ net702 net1018 VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__nand2_1
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20359_ net794 net57 VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__and2_1
XFILLER_136_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11092_ _02034_ _02035_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__nand2_1
XFILLER_95_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14920_ _05818_ _05702_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__nand2_2
XFILLER_102_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14851_ _05670_ _05744_ _05745_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__nand3_2
XFILLER_36_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17570_ _08331_ _08301_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__nand2_1
XFILLER_75_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13802_ net757 net752 net689 net683 VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__and4_1
X_11994_ _02928_ _02858_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__nand2_2
X_16521_ _06878_ _07392_ _07390_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__o21a_1
XFILLER_56_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14782_ net750 net649 VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__nand2_1
X_10945_ net702 net1106 _01889_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__a22o_1
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13733_ _04637_ _04633_ _04630_ _04638_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__o211ai_4
X_16452_ net812 net928 net491 VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__nand3_2
X_10876_ _09690_ net1153 VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__and2_1
XFILLER_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13664_ _04552_ _04567_ _04566_ _04569_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__o211ai_4
X_19240_ _10007_ _10138_ _10139_ VGND VGND VPWR VPWR _10140_ sky130_fd_sc_hd__nand3_4
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16383_ _07226_ _07252_ _07253_ VGND VGND VPWR VPWR _07257_ sky130_fd_sc_hd__nand3_2
X_12615_ _03384_ _03389_ _03386_ VGND VGND VPWR VPWR _03546_ sky130_fd_sc_hd__a21oi_1
X_15403_ _06251_ _06290_ _06295_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__o21bai_2
XTAP_TAPCELL_ROW_14_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19171_ _10030_ _10031_ _10058_ _10059_ VGND VGND VPWR VPWR _10065_ sky130_fd_sc_hd__nand4_2
X_18122_ net790 net781 net601 VGND VGND VPWR VPWR _08970_ sky130_fd_sc_hd__nand3_4
X_13595_ _04409_ _04428_ _04426_ _04424_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__o2bb2ai_2
X_15334_ net730 net912 VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__nand2_1
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12546_ _03463_ _03464_ _03476_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__a21oi_1
XFILLER_61_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18053_ _08876_ _08867_ _08875_ _08864_ _08863_ VGND VGND VPWR VPWR _08902_ sky130_fd_sc_hd__a32o_1
X_12477_ _03396_ _03404_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__nand2_1
X_15265_ net730 net643 VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__and2_1
XANTENNA_4 _00061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ _07868_ _07869_ _07870_ VGND VGND VPWR VPWR _07874_ sky130_fd_sc_hd__a21oi_1
XFILLER_99_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11428_ _09526_ _02363_ net536 net664 _02361_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__o2111ai_4
X_14216_ net676 net670 net1125 _05010_ _05013_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__a32o_2
X_15196_ net733 net909 VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__nand2_1
X_11359_ _02156_ _02292_ _02299_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__o21ai_1
X_14147_ net731 net699 VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__nand2_1
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18955_ _09769_ _09770_ _09844_ _09845_ VGND VGND VPWR VPWR _09847_ sky130_fd_sc_hd__nand4_1
X_14078_ net788 net639 VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__nand2_1
X_17906_ _08727_ _08763_ _08762_ VGND VGND VPWR VPWR _08765_ sky130_fd_sc_hd__a21oi_1
X_13029_ _03944_ _03947_ _03948_ net902 _03954_ VGND VGND VPWR VPWR _03956_ sky130_fd_sc_hd__o2111ai_1
X_18886_ net760 net942 VGND VGND VPWR VPWR _09778_ sky130_fd_sc_hd__nand2_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17837_ net900 net473 _08691_ _08693_ _08687_ VGND VGND VPWR VPWR _08698_ sky130_fd_sc_hd__a41oi_2
XFILLER_67_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer16 net812 VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__buf_1
XFILLER_94_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer27 net823 VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__buf_2
Xrebuffer49 _07507_ VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd1_1
X_17768_ net566 net1054 net484 net480 VGND VGND VPWR VPWR _08630_ sky130_fd_sc_hd__nand4_2
XFILLER_54_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer38 b_l\[9\] VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__buf_4
X_16719_ _07491_ _07549_ _07551_ _07489_ VGND VGND VPWR VPWR _07590_ sky130_fd_sc_hd__a31oi_2
X_17699_ _08558_ _08560_ VGND VGND VPWR VPWR _08562_ sky130_fd_sc_hd__nand2_2
X_19507_ net183 _00588_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__nand2_2
X_19438_ _00620_ _00616_ _00619_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__a21oi_1
X_19369_ net230 VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer106 b_h\[1\] VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__buf_8
Xrebuffer128 _09612_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer117 net912 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer139 a_l\[15\] VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold510 mid_sum\[17\] VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap262 _06748_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_1
Xhold532 p_ll_pipe\[9\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 p_hh\[29\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap240 net241 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
X_20213_ _01451_ _01455_ net794 VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__o21ai_1
Xmax_cap251 _01381_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_1
Xhold554 _00784_ VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 mid_sum\[15\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 term_high\[57\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold576 p_hl\[31\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap284 _06179_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_6
Xmax_cap295 _01144_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_20144_ _09319_ _09351_ _01205_ _01288_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__o31a_1
XFILLER_106_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_20075_ _01299_ _01302_ _01303_ _01222_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10730_ _01760_ _01761_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_45_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10661_ _09537_ _09548_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__nor2_1
XFILLER_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12400_ _03194_ _03197_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10592_ net795 net1309 VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__and2_1
X_13380_ _04286_ _04288_ _04283_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__a21o_1
X_12331_ net1019 b_h\[8\] _03260_ _03263_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a22o_1
X_12262_ _03194_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__nand2_1
X_15050_ _05944_ net677 net719 _05943_ VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__nand4_2
XFILLER_147_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11213_ net691 net517 VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__nand2_1
X_14001_ _04904_ _04906_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__nand2_1
X_12193_ _03006_ _03009_ _03010_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a21oi_1
X_11144_ _02081_ _02083_ _02078_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__a21o_1
XFILLER_96_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput74 net74 VGND VGND VPWR VPWR p[17] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_56_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput85 net85 VGND VGND VPWR VPWR p[27] sky130_fd_sc_hd__buf_2
Xoutput96 net96 VGND VGND VPWR VPWR p[37] sky130_fd_sc_hd__buf_2
X_15952_ _06745_ _06747_ net261 _06821_ _06823_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__o221ai_2
XFILLER_122_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11075_ net702 net517 VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__nand2_1
X_18740_ _09463_ _09594_ _09620_ net300 VGND VGND VPWR VPWR _09627_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18671_ _09547_ _09550_ _09551_ VGND VGND VPWR VPWR _09552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14903_ _05796_ _05799_ _09264_ _09504_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__o2bb2ai_1
X_17622_ _02589_ _07234_ net581 net476 _08484_ VGND VGND VPWR VPWR _08486_ sky130_fd_sc_hd__o2111ai_4
X_15883_ net598 net591 VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__nand2_8
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14834_ _05580_ _05584_ _05730_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__o21ai_4
XFILLER_17_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ net323 _02907_ _02891_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__nand3_1
X_17553_ _08316_ _08325_ _08313_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__o21ai_2
X_14765_ _05663_ _05664_ _05660_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__a21o_1
X_10928_ _01867_ _01873_ _01874_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__nand3b_1
X_16504_ net561 net529 VGND VGND VPWR VPWR _07377_ sky130_fd_sc_hd__nand2_1
X_17484_ _08348_ _08349_ VGND VGND VPWR VPWR _08350_ sky130_fd_sc_hd__nor2_4
X_13716_ _04621_ _04588_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nand2_1
X_16435_ _07180_ _07184_ _07307_ _07308_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__o31a_2
X_19223_ net1128 net717 VGND VGND VPWR VPWR _10121_ sky130_fd_sc_hd__nand2_1
X_14696_ _05595_ _05593_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__nor2_1
X_10859_ net793 net1284 VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__and2_1
X_13647_ net714 net963 _04554_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__and3_1
X_16366_ _07228_ _07238_ _07239_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__nand3_2
X_13578_ _04456_ _04434_ _04435_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__a21oi_4
X_19154_ net765 net568 _10044_ _10045_ VGND VGND VPWR VPWR _10046_ sky130_fd_sc_hd__a22oi_2
XFILLER_145_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16297_ _07168_ _07170_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__nand2_1
X_12529_ _03415_ _03417_ _03457_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__nand3_2
X_18105_ _08936_ _08937_ _08903_ _08899_ VGND VGND VPWR VPWR _08953_ sky130_fd_sc_hd__a31oi_2
X_19085_ _09870_ _09974_ _09975_ VGND VGND VPWR VPWR _09976_ sky130_fd_sc_hd__nand3_4
X_15317_ _06073_ _06146_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__nor2_2
X_18036_ _08884_ _08857_ VGND VGND VPWR VPWR _08886_ sky130_fd_sc_hd__nand2_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15248_ _06079_ _06142_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__nand3b_1
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15179_ _05888_ _05889_ _06075_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__a21boi_1
XFILLER_141_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_19987_ net580 net721 _01208_ _01210_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__a22oi_2
X_18938_ _09827_ _09807_ VGND VGND VPWR VPWR _09830_ sky130_fd_sc_hd__nand2_1
.ends

